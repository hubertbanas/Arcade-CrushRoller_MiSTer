library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"23",X"31",X"B0",X"4F",X"ED",X"56",X"18",X"79",X"A0",X"C3",X"06",X"A0",X"C3",X"09",X"A0",X"C3",
		X"0F",X"0F",X"0F",X"0F",X"C9",X"C3",X"12",X"A0",X"E1",X"D1",X"C1",X"00",X"00",X"C7",X"C3",X"1E",
		X"A0",X"00",X"00",X"00",X"00",X"32",X"3C",X"00",X"00",X"10",X"48",X"00",X"00",X"00",X"00",X"03",
		X"E1",X"22",X"5A",X"4C",X"C9",X"00",X"00",X"18",X"F5",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",
		X"D9",X"C5",X"D5",X"E5",X"08",X"F5",X"21",X"00",X"50",X"36",X"00",X"32",X"C0",X"50",X"2E",X"07",
		X"36",X"01",X"CD",X"D2",X"0B",X"CD",X"DD",X"2B",X"CD",X"D6",X"13",X"CD",X"F7",X"2D",X"CD",X"00",
		X"28",X"CD",X"0D",X"32",X"CD",X"50",X"10",X"3E",X"FF",X"32",X"22",X"4C",X"21",X"00",X"50",X"36",
		X"01",X"F1",X"08",X"E1",X"D1",X"C1",X"D9",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"F1",X"FB",
		X"C9",X"21",X"07",X"50",X"36",X"00",X"2B",X"7C",X"FE",X"3F",X"32",X"C0",X"50",X"20",X"F5",X"16",
		X"00",X"D9",X"21",X"00",X"40",X"36",X"00",X"23",X"7C",X"32",X"C0",X"50",X"FE",X"51",X"20",X"F5",
		X"3E",X"00",X"32",X"03",X"50",X"21",X"00",X"40",X"55",X"5D",X"DD",X"21",X"B1",X"00",X"C3",X"10",
		X"01",X"21",X"00",X"44",X"DD",X"21",X"BB",X"00",X"C3",X"10",X"01",X"21",X"00",X"4C",X"DD",X"21",
		X"C5",X"00",X"C3",X"10",X"01",X"21",X"00",X"40",X"36",X"40",X"23",X"7C",X"FE",X"44",X"20",X"F8",
		X"36",X"03",X"23",X"7C",X"FE",X"48",X"20",X"F8",X"7A",X"B3",X"CA",X"6C",X"01",X"01",X"E0",X"FF",
		X"21",X"A6",X"42",X"36",X"42",X"09",X"36",X"41",X"09",X"36",X"44",X"09",X"36",X"40",X"09",X"36",
		X"52",X"09",X"36",X"41",X"09",X"36",X"4D",X"09",X"36",X"40",X"DD",X"21",X"01",X"01",X"C3",X"4F",
		X"01",X"09",X"53",X"DD",X"21",X"0A",X"01",X"C3",X"4F",X"01",X"16",X"FF",X"D9",X"C3",X"6C",X"01",
		X"7E",X"B7",X"FD",X"21",X"18",X"01",X"20",X"2E",X"3E",X"01",X"47",X"77",X"AE",X"FD",X"21",X"23",
		X"01",X"20",X"23",X"78",X"37",X"8F",X"32",X"C0",X"50",X"30",X"EF",X"23",X"7D",X"06",X"4F",X"32",
		X"07",X"50",X"10",X"FB",X"B7",X"20",X"D9",X"7C",X"FE",X"44",X"28",X"08",X"FE",X"48",X"28",X"04",
		X"FE",X"50",X"20",X"CC",X"DD",X"E9",X"B3",X"5F",X"7A",X"B7",X"20",X"01",X"54",X"FD",X"E9",X"09",
		X"7A",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"37",X"77",X"09",X"7A",
		X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"37",X"77",X"09",X"DD",X"E9",X"21",X"00",X"00",X"11",
		X"04",X"01",X"01",X"00",X"10",X"3E",X"FF",X"AE",X"32",X"07",X"50",X"32",X"C0",X"50",X"23",X"0D",
		X"20",X"F5",X"10",X"F3",X"B7",X"FD",X"21",X"8B",X"01",X"20",X"5A",X"14",X"1D",X"20",X"E3",X"CB",
		X"7A",X"20",X"08",X"D9",X"7A",X"B7",X"20",X"03",X"C3",X"27",X"02",X"21",X"00",X"20",X"10",X"FE",
		X"32",X"C0",X"50",X"2D",X"20",X"F8",X"D9",X"21",X"BA",X"42",X"01",X"E0",X"FF",X"36",X"44",X"09",
		X"36",X"49",X"09",X"36",X"50",X"09",X"09",X"36",X"53",X"09",X"36",X"57",X"09",X"3A",X"00",X"50",
		X"57",X"DD",X"21",X"C8",X"01",X"C3",X"4F",X"01",X"3A",X"40",X"50",X"57",X"DD",X"21",X"D2",X"01",
		X"18",X"F3",X"3A",X"80",X"50",X"57",X"DD",X"21",X"DC",X"01",X"18",X"E9",X"D9",X"25",X"20",X"BE",
		X"C7",X"25",X"20",X"BA",X"C7",X"08",X"7A",X"87",X"CB",X"FA",X"E6",X"3F",X"D9",X"21",X"A8",X"42",
		X"85",X"6F",X"30",X"01",X"24",X"01",X"E0",X"FF",X"36",X"42",X"09",X"36",X"41",X"09",X"36",X"44",
		X"09",X"09",X"36",X"50",X"09",X"36",X"52",X"09",X"36",X"4F",X"09",X"36",X"4D",X"09",X"D9",X"7A",
		X"D9",X"E6",X"0F",X"57",X"DD",X"21",X"1B",X"02",X"C3",X"4F",X"01",X"08",X"57",X"DD",X"21",X"24",
		X"02",X"C3",X"4F",X"01",X"D9",X"FD",X"E9",X"CD",X"D7",X"2D",X"CD",X"03",X"38",X"CD",X"00",X"38",
		X"CD",X"66",X"0B",X"21",X"00",X"10",X"06",X"2F",X"7D",X"32",X"C0",X"50",X"32",X"07",X"50",X"10",
		X"F7",X"2B",X"7D",X"B4",X"20",X"F0",X"21",X"00",X"40",X"36",X"00",X"23",X"7C",X"FE",X"51",X"20",
		X"F8",X"3E",X"03",X"CD",X"5B",X"2E",X"3E",X"40",X"CD",X"65",X"2E",X"3E",X"01",X"32",X"00",X"50",
		X"3A",X"80",X"50",X"32",X"00",X"4C",X"CD",X"E7",X"1B",X"CD",X"2A",X"2E",X"3E",X"08",X"32",X"20",
		X"4C",X"CD",X"A8",X"1D",X"CD",X"9F",X"1C",X"FB",X"CD",X"D7",X"2D",X"21",X"90",X"4C",X"CD",X"5F",
		X"39",X"7E",X"35",X"B7",X"20",X"5C",X"34",X"21",X"20",X"4C",X"3A",X"1E",X"4C",X"B7",X"28",X"0B",
		X"7E",X"E6",X"03",X"20",X"06",X"CC",X"54",X"0C",X"C3",X"86",X"03",X"AF",X"32",X"AD",X"4C",X"CB",
		X"7E",X"C4",X"9F",X"03",X"21",X"20",X"4C",X"7E",X"CB",X"77",X"E5",X"C4",X"7F",X"04",X"E1",X"CB",
		X"6E",X"E5",X"C4",X"24",X"04",X"E1",X"7E",X"E6",X"03",X"20",X"11",X"CB",X"5E",X"28",X"0D",X"3A",
		X"AC",X"4C",X"B7",X"00",X"00",X"00",X"CD",X"75",X"05",X"F2",X"89",X"03",X"21",X"87",X"4C",X"7E",
		X"35",X"B7",X"20",X"35",X"3A",X"5C",X"4C",X"FE",X"01",X"20",X"04",X"36",X"01",X"18",X"2A",X"34",
		X"18",X"29",X"21",X"C4",X"4F",X"47",X"FE",X"FF",X"20",X"02",X"36",X"CC",X"E6",X"9F",X"FE",X"9F",
		X"20",X"05",X"7E",X"C6",X"04",X"18",X"0F",X"78",X"E6",X"1F",X"FE",X"1F",X"20",X"7F",X"CB",X"68",
		X"3E",X"DC",X"28",X"02",X"3E",X"78",X"77",X"18",X"74",X"18",X"7E",X"CD",X"52",X"1D",X"3A",X"80",
		X"50",X"CB",X"6F",X"20",X"06",X"CD",X"4A",X"3B",X"CD",X"17",X"3C",X"CD",X"55",X"2D",X"CD",X"4F",
		X"0A",X"CD",X"E1",X"08",X"CD",X"8F",X"08",X"CD",X"B7",X"08",X"CD",X"1B",X"18",X"CD",X"00",X"08",
		X"3A",X"06",X"4E",X"FE",X"01",X"D4",X"E0",X"1A",X"CD",X"AA",X"0D",X"CD",X"5B",X"1C",X"CD",X"3F",
		X"24",X"CD",X"C6",X"15",X"CD",X"86",X"39",X"CD",X"40",X"26",X"CD",X"B0",X"1B",X"CD",X"27",X"13",
		X"CD",X"AA",X"14",X"CD",X"1D",X"0A",X"CD",X"81",X"09",X"CD",X"F1",X"3A",X"CD",X"93",X"2A",X"CD",
		X"06",X"38",X"CD",X"7D",X"12",X"CD",X"CC",X"10",X"CD",X"75",X"10",X"CD",X"6A",X"11",X"CD",X"0A",
		X"20",X"CD",X"6C",X"23",X"CD",X"B6",X"1C",X"CD",X"C0",X"19",X"CD",X"E4",X"2A",X"CD",X"97",X"2C",
		X"CD",X"ED",X"2C",X"CD",X"F6",X"11",X"CD",X"BC",X"23",X"CD",X"FC",X"23",X"CD",X"4C",X"2E",X"AF",
		X"32",X"22",X"4C",X"3A",X"22",X"4C",X"B7",X"32",X"C0",X"50",X"C2",X"7B",X"02",X"18",X"F4",X"3E",
		X"43",X"CD",X"5B",X"2E",X"AF",X"32",X"A2",X"4C",X"CD",X"2A",X"2E",X"21",X"B0",X"4F",X"06",X"50",
		X"CD",X"C5",X"2D",X"21",X"80",X"4E",X"CD",X"C5",X"2D",X"32",X"8E",X"4C",X"CD",X"6F",X"2E",X"CD",
		X"00",X"10",X"CD",X"5A",X"2C",X"3E",X"80",X"32",X"CE",X"4F",X"21",X"00",X"4E",X"06",X"40",X"CD",
		X"C5",X"2D",X"CD",X"38",X"22",X"3E",X"05",X"32",X"0E",X"4E",X"21",X"20",X"4C",X"7E",X"E6",X"03",
		X"CB",X"BE",X"CA",X"1B",X"24",X"CD",X"B1",X"2D",X"CD",X"B9",X"2D",X"3E",X"C0",X"32",X"87",X"4C",
		X"21",X"10",X"40",X"06",X"10",X"CD",X"66",X"23",X"CD",X"AC",X"21",X"CD",X"EA",X"39",X"CD",X"38",
		X"22",X"3E",X"81",X"32",X"5C",X"4C",X"3E",X"C7",X"32",X"AE",X"4C",X"CD",X"D7",X"2D",X"3A",X"C0",
		X"50",X"E6",X"30",X"FE",X"10",X"C9",X"3A",X"80",X"50",X"E6",X"C0",X"C8",X"00",X"00",X"21",X"12",
		X"4E",X"36",X"30",X"C9",X"CB",X"AE",X"E5",X"CD",X"C6",X"12",X"21",X"B0",X"4F",X"06",X"50",X"CD",
		X"C5",X"2D",X"CD",X"42",X"2F",X"CD",X"6F",X"2E",X"CD",X"00",X"10",X"CD",X"5A",X"2C",X"21",X"03",
		X"4E",X"06",X"03",X"CD",X"C5",X"2D",X"34",X"23",X"77",X"23",X"77",X"32",X"10",X"4E",X"32",X"11",
		X"4E",X"32",X"1B",X"4E",X"3E",X"C0",X"32",X"87",X"4C",X"CD",X"EA",X"39",X"CD",X"38",X"22",X"CD",
		X"9D",X"23",X"CD",X"AC",X"21",X"01",X"3F",X"C0",X"3E",X"80",X"32",X"CE",X"4F",X"E1",X"3A",X"C1",
		X"50",X"A1",X"B9",X"C9",X"3A",X"80",X"50",X"A0",X"B8",X"C8",X"00",X"00",X"C3",X"C3",X"2B",X"CB",
		X"B6",X"E5",X"4E",X"3E",X"03",X"A1",X"28",X"56",X"EB",X"21",X"B0",X"4F",X"06",X"50",X"CD",X"C5",
		X"2D",X"21",X"07",X"4E",X"7E",X"B7",X"28",X"12",X"E6",X"81",X"EA",X"AA",X"04",X"3A",X"12",X"4E",
		X"FE",X"20",X"30",X"04",X"36",X"00",X"18",X"02",X"36",X"FF",X"21",X"1C",X"4C",X"CB",X"51",X"20",
		X"16",X"35",X"20",X"0D",X"CB",X"81",X"CB",X"49",X"20",X"3C",X"C5",X"CD",X"B1",X"2D",X"C1",X"18",
		X"1D",X"CB",X"49",X"20",X"31",X"18",X"62",X"23",X"35",X"20",X"0D",X"CB",X"89",X"CB",X"41",X"20",
		X"36",X"C5",X"CD",X"B9",X"2D",X"C1",X"18",X"06",X"CB",X"41",X"20",X"2B",X"18",X"4B",X"CD",X"E0",
		X"2D",X"3E",X"00",X"32",X"5C",X"4C",X"CB",X"D9",X"CB",X"91",X"CD",X"D7",X"2D",X"E1",X"71",X"3E",
		X"81",X"32",X"AC",X"4C",X"18",X"52",X"E5",X"D5",X"C5",X"CD",X"E5",X"3B",X"CD",X"F1",X"25",X"CD",
		X"B1",X"2D",X"CD",X"A9",X"2D",X"18",X"0F",X"E5",X"D5",X"C5",X"CD",X"E5",X"3B",X"CD",X"F1",X"25",
		X"CD",X"B9",X"2D",X"CD",X"A1",X"2D",X"C1",X"D1",X"E1",X"3E",X"04",X"A9",X"EB",X"77",X"CD",X"6C",
		X"24",X"CD",X"27",X"26",X"CD",X"61",X"3C",X"18",X"02",X"EB",X"71",X"CD",X"5A",X"2C",X"E1",X"3A",
		X"00",X"50",X"CB",X"67",X"20",X"05",X"CD",X"D7",X"2D",X"18",X"08",X"CB",X"56",X"CC",X"D7",X"2D",
		X"C4",X"DA",X"2D",X"3E",X"81",X"32",X"5C",X"4C",X"3E",X"8F",X"32",X"87",X"4C",X"CD",X"EA",X"39",
		X"CD",X"38",X"22",X"CD",X"AC",X"21",X"CD",X"29",X"10",X"3E",X"80",X"32",X"CE",X"4F",X"0E",X"C0",
		X"3A",X"C2",X"50",X"E6",X"3F",X"FE",X"2F",X"C9",X"3A",X"81",X"50",X"A1",X"B9",X"C0",X"00",X"00",
		X"21",X"03",X"4E",X"35",X"C9",X"CD",X"C5",X"05",X"21",X"87",X"4C",X"36",X"C0",X"21",X"C0",X"4F",
		X"7E",X"B7",X"20",X"06",X"CD",X"50",X"0D",X"C3",X"E1",X"05",X"FE",X"01",X"CA",X"05",X"06",X"FE",
		X"03",X"CA",X"5D",X"06",X"FE",X"07",X"CA",X"09",X"38",X"FE",X"0F",X"CA",X"51",X"39",X"FE",X"1F",
		X"C0",X"3E",X"80",X"32",X"20",X"4C",X"AF",X"32",X"C0",X"4F",X"32",X"A2",X"4C",X"32",X"C1",X"4F",
		X"3A",X"C3",X"50",X"E6",X"3F",X"FE",X"3C",X"C9",X"3A",X"85",X"50",X"E6",X"C0",X"FE",X"C0",X"C8",
		X"00",X"00",X"C2",X"5D",X"06",X"21",X"A2",X"4C",X"7E",X"FE",X"0A",X"D0",X"3A",X"83",X"4C",X"E6",
		X"1F",X"FE",X"10",X"C0",X"7E",X"34",X"FE",X"04",X"CA",X"DF",X"0C",X"FE",X"06",X"CA",X"02",X"0D",
		X"C9",X"21",X"C4",X"4F",X"36",X"FA",X"23",X"36",X"01",X"21",X"E4",X"4F",X"36",X"FF",X"23",X"36",
		X"CC",X"3E",X"81",X"32",X"CE",X"4F",X"3E",X"01",X"32",X"C0",X"4F",X"3E",X"06",X"32",X"19",X"4E",
		X"AF",X"32",X"06",X"4E",X"C9",X"21",X"D4",X"4F",X"36",X"44",X"CD",X"40",X"26",X"CD",X"E4",X"2A",
		X"21",X"E4",X"4F",X"7E",X"FE",X"02",X"30",X"06",X"3E",X"03",X"32",X"C0",X"4F",X"C9",X"E6",X"06",
		X"C0",X"7E",X"E6",X"FE",X"21",X"47",X"06",X"06",X"0B",X"BE",X"23",X"28",X"04",X"23",X"10",X"F9",
		X"C9",X"7E",X"F5",X"21",X"E4",X"4F",X"CD",X"7F",X"2C",X"21",X"00",X"40",X"19",X"F1",X"2B",X"77",
		X"7C",X"C6",X"04",X"67",X"36",X"01",X"C9",X"B8",X"43",X"B0",X"52",X"A8",X"55",X"A0",X"53",X"98",
		X"48",X"88",X"52",X"80",X"4F",X"78",X"4C",X"70",X"4C",X"68",X"45",X"60",X"52",X"01",X"F8",X"1C",
		X"21",X"53",X"40",X"CD",X"9F",X"06",X"0E",X"FF",X"23",X"CD",X"9F",X"06",X"23",X"CD",X"9F",X"06",
		X"0E",X"F7",X"23",X"CD",X"9F",X"06",X"21",X"73",X"41",X"01",X"5B",X"0A",X"CD",X"9F",X"06",X"21",
		X"76",X"41",X"0E",X"EE",X"CD",X"9F",X"06",X"21",X"54",X"40",X"36",X"D2",X"23",X"36",X"FC",X"21",
		X"B4",X"43",X"36",X"FE",X"23",X"36",X"FD",X"3E",X"07",X"32",X"C0",X"4F",X"C3",X"DA",X"2E",X"C5",
		X"E5",X"11",X"20",X"00",X"71",X"19",X"10",X"FC",X"E1",X"C1",X"C9",X"CD",X"ED",X"06",X"2A",X"80",
		X"4C",X"E5",X"3A",X"82",X"4C",X"F5",X"CD",X"D2",X"06",X"CD",X"C6",X"12",X"F1",X"32",X"82",X"4C",
		X"E1",X"22",X"80",X"4C",X"CD",X"4C",X"2E",X"C9",X"3A",X"06",X"4E",X"3C",X"FE",X"09",X"D8",X"3E",
		X"09",X"C9",X"CD",X"C8",X"06",X"21",X"80",X"4C",X"36",X"00",X"23",X"77",X"23",X"36",X"00",X"21",
		X"01",X"4E",X"86",X"27",X"77",X"D0",X"2B",X"7E",X"C6",X"01",X"27",X"77",X"C9",X"CD",X"E9",X"2D",
		X"08",X"CC",X"43",X"53",X"55",X"4E",X"4F",X"42",X"40",X"40",X"40",X"C9",X"00",X"00",X"18",X"96",
		X"EB",X"CD",X"E9",X"1A",X"21",X"A8",X"05",X"E3",X"E5",X"EB",X"23",X"0E",X"0A",X"C3",X"C3",X"21",
		X"3A",X"2F",X"02",X"B7",X"28",X"0B",X"CD",X"26",X"15",X"38",X"0D",X"CD",X"20",X"19",X"C3",X"DE",
		X"04",X"CD",X"1F",X"15",X"38",X"09",X"18",X"14",X"2A",X"3E",X"00",X"7C",X"B5",X"20",X"0D",X"2A",
		X"40",X"00",X"7C",X"B5",X"28",X"22",X"CD",X"59",X"18",X"C3",X"FE",X"1B",X"7E",X"23",X"5E",X"16",
		X"00",X"23",X"E5",X"21",X"9B",X"22",X"19",X"19",X"5E",X"23",X"56",X"EB",X"E3",X"CB",X"67",X"C8",
		X"3A",X"52",X"00",X"B7",X"C8",X"C3",X"21",X"1B",X"06",X"04",X"AF",X"CD",X"61",X"1B",X"10",X"FB",
		X"3E",X"4F",X"CD",X"30",X"1B",X"C3",X"1E",X"12",X"CD",X"AE",X"18",X"F5",X"C5",X"CD",X"E5",X"16",
		X"38",X"07",X"CD",X"66",X"18",X"38",X"11",X"B6",X"57",X"C1",X"F1",X"38",X"12",X"B2",X"57",X"FE",
		X"76",X"CC",X"01",X"1B",X"7A",X"C3",X"61",X"1B",X"B6",X"57",X"F1",X"F1",X"DC",X"01",X"1B",X"B2",
		X"57",X"FE",X"76",X"CC",X"01",X"1B",X"78",X"CD",X"61",X"1B",X"7A",X"CD",X"61",X"1B",X"79",X"C3",
		X"61",X"1B",X"CD",X"AE",X"18",X"38",X"0D",X"B6",X"CD",X"61",X"1B",X"CD",X"BB",X"16",X"CD",X"0C",
		X"19",X"C3",X"61",X"1B",X"B6",X"CD",X"90",X"07",X"18",X"F1",X"CD",X"AE",X"18",X"38",X"04",X"B6",
		X"C3",X"61",X"1B",X"B6",X"C3",X"90",X"07",X"CD",X"66",X"18",X"18",X"F1",X"7E",X"C3",X"61",X"1B",
		X"7E",X"CD",X"61",X"1B",X"23",X"18",X"F5",X"7E",X"CD",X"61",X"1B",X"CD",X"A4",X"14",X"18",X"CE",
		X"CD",X"F7",X"18",X"B6",X"CD",X"61",X"1B",X"CD",X"BB",X"16",X"CD",X"98",X"1E",X"C3",X"FE",X"1B",
		X"7E",X"CD",X"61",X"1B",X"CD",X"A4",X"14",X"18",X"F1",X"CD",X"CF",X"18",X"30",X"E5",X"57",X"24",
		X"21",X"E4",X"4F",X"7E",X"FE",X"88",X"28",X"09",X"23",X"7E",X"FE",X"60",X"28",X"03",X"FE",X"C0",
		X"C0",X"21",X"E8",X"4F",X"CD",X"1A",X"08",X"21",X"EA",X"4F",X"E5",X"CD",X"6B",X"08",X"E1",X"79",
		X"B7",X"C8",X"7D",X"D6",X"10",X"6F",X"3A",X"1B",X"4E",X"FE",X"02",X"38",X"24",X"FE",X"04",X"38",
		X"0D",X"E5",X"7D",X"C6",X"10",X"6F",X"7E",X"23",X"B6",X"E6",X"07",X"E1",X"28",X"18",X"E5",X"7D",
		X"C6",X"10",X"6F",X"7E",X"FE",X"88",X"20",X"02",X"23",X"7E",X"E6",X"0F",X"FE",X"08",X"E1",X"28",
		X"05",X"7E",X"CD",X"FE",X"18",X"C8",X"3A",X"11",X"4E",X"B7",X"F5",X"C4",X"FD",X"3A",X"F1",X"CC",
		X"73",X"0D",X"7E",X"D7",X"E6",X"0F",X"A1",X"C8",X"23",X"71",X"C9",X"11",X"E4",X"4F",X"0E",X"00",
		X"1A",X"BE",X"28",X"10",X"23",X"13",X"1A",X"BE",X"C0",X"2B",X"1B",X"1A",X"96",X"07",X"0E",X"04",
		X"D8",X"0E",X"02",X"C9",X"23",X"13",X"1A",X"96",X"07",X"0E",X"08",X"D8",X"0E",X"01",X"C9",X"21",
		X"E8",X"4F",X"CD",X"BE",X"1A",X"20",X"1B",X"E5",X"7D",X"D6",X"10",X"6F",X"7E",X"E6",X"F0",X"5F",
		X"D7",X"57",X"7E",X"E6",X"0F",X"20",X"0A",X"ED",X"5F",X"CD",X"58",X"10",X"79",X"A2",X"B3",X"23",
		X"77",X"E1",X"CD",X"48",X"2D",X"18",X"DB",X"3A",X"20",X"4C",X"E6",X"07",X"C0",X"21",X"D4",X"4F",
		X"7E",X"CD",X"FE",X"18",X"C8",X"7E",X"CD",X"CC",X"08",X"23",X"77",X"C9",X"E6",X"06",X"0E",X"06",
		X"28",X"02",X"0E",X"09",X"ED",X"5F",X"0F",X"0F",X"06",X"0C",X"38",X"02",X"06",X"03",X"79",X"A0",
		X"C9",X"21",X"EC",X"4F",X"CD",X"BE",X"1A",X"C0",X"56",X"23",X"5E",X"21",X"08",X"09",X"01",X"FF",
		X"09",X"7E",X"BA",X"23",X"20",X"02",X"7E",X"BB",X"23",X"28",X"05",X"23",X"10",X"F3",X"18",X"01",
		X"4E",X"21",X"DC",X"4F",X"7E",X"A1",X"77",X"C9",X"88",X"D8",X"7F",X"58",X"C0",X"DF",X"B8",X"C0",
		X"BF",X"68",X"98",X"CF",X"B8",X"98",X"BF",X"88",X"78",X"6F",X"58",X"60",X"CF",X"B8",X"60",X"3F",
		X"88",X"38",X"EF",X"21",X"E4",X"4F",X"7E",X"FE",X"88",X"23",X"20",X"0B",X"7E",X"2B",X"FE",X"80",
		X"28",X"14",X"FE",X"D0",X"C0",X"18",X"19",X"7E",X"FE",X"60",X"C0",X"2B",X"7E",X"FE",X"60",X"28",
		X"19",X"FE",X"B0",X"C0",X"18",X"1E",X"01",X"BD",X"11",X"11",X"88",X"80",X"21",X"F0",X"41",X"C9",
		X"01",X"BC",X"18",X"11",X"88",X"D0",X"21",X"E7",X"41",X"C9",X"01",X"BA",X"12",X"11",X"60",X"60",
		X"21",X"74",X"41",X"C9",X"01",X"B8",X"14",X"11",X"B0",X"60",X"21",X"94",X"42",X"3A",X"4F",X"50",
		X"07",X"C9",X"3A",X"90",X"50",X"E6",X"C0",X"C8",X"87",X"87",X"D8",X"00",X"00",X"21",X"34",X"42",
		X"C9",X"3A",X"40",X"50",X"0F",X"38",X"12",X"3A",X"83",X"4C",X"FE",X"4F",X"20",X"0B",X"CD",X"D0",
		X"3A",X"28",X"06",X"00",X"00",X"32",X"03",X"4E",X"E5",X"3A",X"11",X"4E",X"B7",X"C8",X"21",X"E6",
		X"4F",X"CD",X"3F",X"2C",X"CD",X"BE",X"1A",X"28",X"07",X"3A",X"83",X"4C",X"0F",X"DC",X"3F",X"2C",
		X"E5",X"E5",X"E5",X"CD",X"FF",X"09",X"E1",X"11",X"E4",X"4F",X"01",X"02",X"00",X"ED",X"B0",X"3A",
		X"D6",X"4F",X"32",X"D4",X"4F",X"E1",X"CD",X"26",X"09",X"28",X"02",X"E1",X"C9",X"78",X"0F",X"F5",
		X"DC",X"F2",X"2E",X"F1",X"0F",X"F5",X"DC",X"E2",X"2E",X"F1",X"0F",X"F5",X"DC",X"DA",X"2E",X"F1",
		X"0F",X"DC",X"FA",X"2E",X"E1",X"AF",X"77",X"23",X"77",X"32",X"C6",X"4F",X"32",X"D6",X"4F",X"32",
		X"11",X"4E",X"E5",X"CD",X"D1",X"31",X"21",X"9D",X"4C",X"36",X"FF",X"23",X"34",X"E1",X"C9",X"3A",
		X"83",X"4C",X"21",X"C6",X"4F",X"CB",X"56",X"28",X"0A",X"CB",X"57",X"28",X"03",X"CB",X"8E",X"C9",
		X"CB",X"CE",X"C9",X"CB",X"57",X"28",X"03",X"CB",X"86",X"C9",X"CB",X"C6",X"C9",X"CD",X"23",X"09",
		X"C0",X"7E",X"CD",X"B2",X"16",X"D0",X"3A",X"D4",X"4F",X"E6",X"0F",X"A0",X"C8",X"78",X"32",X"D6",
		X"4F",X"79",X"32",X"11",X"4E",X"32",X"C6",X"4F",X"3E",X"03",X"32",X"C7",X"4F",X"E5",X"CD",X"C9",
		X"31",X"E1",X"ED",X"53",X"E6",X"4F",X"78",X"E6",X"06",X"CA",X"2E",X"2F",X"C3",X"28",X"2F",X"21",
		X"E4",X"4F",X"CD",X"BE",X"1A",X"20",X"38",X"DD",X"21",X"00",X"40",X"CD",X"7F",X"2C",X"FD",X"21",
		X"00",X"44",X"DD",X"19",X"FD",X"19",X"0E",X"00",X"CD",X"94",X"0A",X"CB",X"09",X"CD",X"B4",X"0A",
		X"CB",X"09",X"CD",X"D4",X"0A",X"CB",X"09",X"CD",X"F4",X"0A",X"CB",X"09",X"CD",X"40",X"0B",X"E5",
		X"7D",X"D6",X"10",X"6F",X"3E",X"0F",X"A6",X"47",X"79",X"D7",X"E6",X"F0",X"B0",X"77",X"E1",X"CD",
		X"48",X"2D",X"18",X"BE",X"FD",X"56",X"FE",X"FD",X"5E",X"1E",X"CD",X"27",X"0B",X"DD",X"56",X"FE",
		X"DD",X"5E",X"1E",X"CD",X"B5",X"22",X"3E",X"D1",X"CD",X"E6",X"22",X"3E",X"EA",X"CD",X"E6",X"22",
		X"CD",X"14",X"0B",X"C9",X"FD",X"56",X"40",X"FD",X"5E",X"3F",X"CD",X"27",X"0B",X"DD",X"56",X"40",
		X"DD",X"5E",X"3F",X"CD",X"B5",X"22",X"3E",X"E1",X"CD",X"E6",X"22",X"3E",X"E5",X"CD",X"E6",X"22",
		X"CD",X"14",X"0B",X"C9",X"FD",X"56",X"E0",X"FD",X"5E",X"DF",X"CD",X"27",X"0B",X"DD",X"56",X"E0",
		X"DD",X"5E",X"DF",X"CD",X"B5",X"22",X"3E",X"E5",X"CD",X"E6",X"22",X"3E",X"E1",X"CD",X"E6",X"22",
		X"CD",X"14",X"0B",X"C9",X"FD",X"56",X"01",X"FD",X"5E",X"21",X"CD",X"27",X"0B",X"DD",X"56",X"01",
		X"DD",X"5E",X"21",X"CD",X"B5",X"22",X"3E",X"EA",X"CD",X"E6",X"22",X"3E",X"D1",X"CD",X"E6",X"22",
		X"CD",X"14",X"0B",X"C9",X"7B",X"FE",X"D8",X"D8",X"FE",X"E0",X"D0",X"7A",X"FE",X"D8",X"D8",X"FE",
		X"E0",X"D0",X"CB",X"E1",X"33",X"33",X"C9",X"7B",X"E6",X"1F",X"FE",X"03",X"28",X"05",X"CD",X"47",
		X"1D",X"20",X"0A",X"7A",X"E6",X"1F",X"FE",X"03",X"C8",X"CD",X"47",X"1D",X"C8",X"33",X"33",X"C9",
		X"06",X"00",X"7E",X"FE",X"88",X"23",X"20",X"0E",X"7E",X"FE",X"10",X"20",X"02",X"CB",X"D8",X"7E",
		X"FE",X"00",X"20",X"02",X"CB",X"C0",X"2B",X"7E",X"FE",X"21",X"38",X"04",X"FE",X"F0",X"38",X"02",
		X"06",X"06",X"78",X"B1",X"4F",X"C9",X"21",X"F0",X"4F",X"06",X"10",X"36",X"00",X"23",X"10",X"FB",
		X"21",X"00",X"40",X"11",X"40",X"F9",X"CD",X"C5",X"0B",X"11",X"F8",X"F2",X"CD",X"C5",X"0B",X"11",
		X"F2",X"F9",X"CD",X"C5",X"0B",X"11",X"F8",X"40",X"CD",X"C5",X"0B",X"7C",X"FE",X"43",X"20",X"EF",
		X"7D",X"FE",X"80",X"20",X"EA",X"11",X"F2",X"F9",X"CD",X"C5",X"0B",X"11",X"F4",X"FA",X"CD",X"C5",
		X"0B",X"11",X"F7",X"F1",X"CD",X"C5",X"0B",X"11",X"F8",X"F2",X"CD",X"C5",X"0B",X"3E",X"F4",X"32",
		X"3D",X"40",X"32",X"FD",X"43",X"3E",X"FA",X"32",X"1D",X"40",X"3E",X"F3",X"32",X"DD",X"43",X"3E",
		X"0B",X"CD",X"5B",X"2E",X"C9",X"72",X"23",X"73",X"23",X"7D",X"E6",X"1F",X"20",X"F7",X"32",X"C0",
		X"50",X"C9",X"CD",X"44",X"0C",X"3A",X"00",X"4C",X"E6",X"03",X"28",X"62",X"3A",X"00",X"50",X"CB",
		X"77",X"21",X"19",X"4C",X"CD",X"F7",X"0B",X"3A",X"00",X"50",X"CB",X"6F",X"21",X"1A",X"4C",X"CD",
		X"F7",X"0B",X"3A",X"00",X"50",X"CB",X"7F",X"7E",X"28",X"05",X"E6",X"0F",X"C8",X"35",X"C9",X"E6",
		X"0F",X"CB",X"D6",X"CB",X"8E",X"C0",X"3A",X"00",X"4C",X"E6",X"03",X"47",X"3A",X"1E",X"4C",X"05",
		X"28",X"0B",X"05",X"28",X"2B",X"7E",X"C6",X"80",X"77",X"D0",X"3A",X"1E",X"4C",X"C6",X"01",X"27",
		X"30",X"02",X"3E",X"99",X"32",X"1E",X"4C",X"3A",X"40",X"50",X"87",X"C9",X"3A",X"80",X"50",X"E6",
		X"C0",X"C8",X"CB",X"77",X"C0",X"00",X"00",X"32",X"19",X"4E",X"32",X"1E",X"4C",X"C9",X"3E",X"97",
		X"C6",X"02",X"18",X"DB",X"21",X"83",X"4C",X"7E",X"FE",X"02",X"D0",X"2F",X"32",X"07",X"50",X"0F",
		X"D8",X"C3",X"B5",X"3A",X"3A",X"AE",X"4C",X"B7",X"18",X"03",X"C3",X"C4",X"1D",X"3A",X"AD",X"4C",
		X"B7",X"20",X"07",X"3C",X"32",X"AD",X"4C",X"C3",X"50",X"0D",X"3A",X"1E",X"4C",X"3D",X"20",X"15",
		X"CD",X"80",X"28",X"0D",X"0F",X"41",X"59",X"4C",X"4E",X"4F",X"40",X"52",X"45",X"59",X"41",X"4C",
		X"50",X"40",X"01",X"18",X"14",X"CD",X"80",X"28",X"0E",X"0F",X"41",X"53",X"52",X"45",X"59",X"41",
		X"4C",X"50",X"40",X"02",X"40",X"52",X"4F",X"40",X"01",X"CD",X"80",X"28",X"11",X"CC",X"40",X"4E",
		X"4F",X"54",X"54",X"55",X"42",X"40",X"54",X"52",X"41",X"54",X"53",X"40",X"48",X"53",X"55",X"50",
		X"CD",X"DF",X"0C",X"CD",X"02",X"0D",X"CD",X"BF",X"0C",X"3E",X"FF",X"32",X"AD",X"4C",X"C9",X"CD",
		X"80",X"28",X"0C",X"47",X"41",X"52",X"45",X"4C",X"4C",X"4F",X"52",X"40",X"48",X"53",X"55",X"52",
		X"43",X"21",X"47",X"45",X"11",X"20",X"00",X"06",X"0C",X"36",X"01",X"19",X"10",X"FB",X"C9",X"CD",
		X"80",X"28",X"09",X"9A",X"41",X"52",X"45",X"56",X"4F",X"40",X"45",X"4D",X"41",X"47",X"21",X"9A",
		X"45",X"01",X"05",X"0F",X"CD",X"9F",X"06",X"21",X"15",X"40",X"06",X"09",X"36",X"40",X"23",X"10",
		X"FB",X"C9",X"CD",X"80",X"28",X"18",X"BC",X"40",X"40",X"44",X"54",X"4C",X"40",X"43",X"49",X"52",
		X"54",X"43",X"45",X"4C",X"45",X"40",X"4F",X"43",X"53",X"45",X"40",X"4C",X"41",X"52",X"55",X"4B",
		X"21",X"BC",X"44",X"01",X"07",X"18",X"CD",X"9F",X"06",X"21",X"E2",X"4F",X"36",X"E8",X"23",X"36",
		X"30",X"21",X"C2",X"4F",X"36",X"04",X"23",X"36",X"07",X"CD",X"80",X"28",X"04",X"FB",X"42",X"01",
		X"08",X"09",X"01",X"21",X"FB",X"46",X"06",X"04",X"36",X"07",X"CD",X"50",X"21",X"10",X"F9",X"C9",
		X"21",X"40",X"40",X"01",X"7F",X"04",X"3E",X"40",X"C5",X"CD",X"D1",X"2D",X"C1",X"3E",X"03",X"21",
		X"40",X"44",X"CD",X"D1",X"2D",X"06",X"50",X"21",X"B0",X"4F",X"CD",X"C5",X"2D",X"CD",X"1B",X"24",
		X"C3",X"38",X"22",X"3A",X"1B",X"4E",X"FE",X"04",X"D8",X"3A",X"06",X"4E",X"B7",X"C8",X"E5",X"7D",
		X"C6",X"11",X"6F",X"7E",X"E1",X"FE",X"60",X"C0",X"3A",X"E5",X"4F",X"FE",X"60",X"C0",X"3A",X"E4",
		X"4F",X"FE",X"58",X"28",X"0C",X"FE",X"B8",X"C0",X"3A",X"94",X"42",X"FE",X"DE",X"C0",X"0E",X"04",
		X"C9",X"3A",X"74",X"41",X"FE",X"DC",X"C0",X"0E",X"02",X"C9",X"3A",X"1B",X"4E",X"FE",X"05",X"D8",
		X"21",X"45",X"0E",X"FE",X"07",X"38",X"0A",X"21",X"6D",X"0E",X"FE",X"09",X"38",X"03",X"21",X"95",
		X"0E",X"D9",X"11",X"E4",X"4F",X"21",X"E8",X"4F",X"D9",X"E5",X"CD",X"D3",X"0D",X"E1",X"D9",X"21",
		X"EA",X"4F",X"D9",X"01",X"00",X"04",X"E5",X"CD",X"F9",X"0D",X"E1",X"79",X"B7",X"20",X"08",X"3E",
		X"0A",X"CD",X"52",X"21",X"10",X"F0",X"C9",X"D9",X"7D",X"D6",X"10",X"6F",X"7E",X"D7",X"E6",X"0F",
		X"D9",X"A1",X"D9",X"28",X"02",X"23",X"77",X"D9",X"C9",X"D9",X"1A",X"96",X"30",X"02",X"ED",X"44",
		X"FE",X"14",X"D9",X"30",X"0F",X"D9",X"23",X"13",X"1A",X"96",X"30",X"02",X"ED",X"44",X"FE",X"14",
		X"2B",X"1B",X"D9",X"D8",X"5E",X"23",X"56",X"23",X"1A",X"BE",X"C0",X"23",X"7E",X"23",X"B7",X"28",
		X"06",X"D9",X"BE",X"D9",X"C0",X"18",X"07",X"7E",X"D9",X"23",X"BE",X"2B",X"D9",X"C0",X"23",X"D9",
		X"1A",X"D9",X"BE",X"D0",X"23",X"BE",X"D8",X"23",X"D9",X"13",X"1A",X"1B",X"D9",X"BE",X"D0",X"23",
		X"BE",X"D8",X"23",X"4E",X"C9",X"94",X"42",X"DE",X"00",X"60",X"B9",X"AF",X"64",X"58",X"04",X"74",
		X"41",X"DC",X"00",X"60",X"69",X"5F",X"68",X"5C",X"02",X"10",X"42",X"DB",X"88",X"00",X"8C",X"84",
		X"80",X"78",X"01",X"07",X"42",X"D9",X"88",X"00",X"8C",X"84",X"D4",X"D0",X"08",X"94",X"42",X"DE",
		X"00",X"60",X"BC",X"AC",X"70",X"58",X"04",X"74",X"41",X"DC",X"00",X"60",X"64",X"57",X"68",X"58",
		X"02",X"10",X"42",X"DB",X"88",X"00",X"94",X"7C",X"84",X"74",X"01",X"07",X"42",X"D9",X"88",X"00",
		X"94",X"7C",X"DC",X"CC",X"08",X"94",X"42",X"DE",X"00",X"60",X"C9",X"9C",X"77",X"58",X"04",X"74",
		X"41",X"DC",X"00",X"60",X"78",X"48",X"68",X"48",X"02",X"10",X"42",X"DB",X"88",X"00",X"A0",X"70",
		X"A0",X"70",X"01",X"07",X"42",X"D9",X"88",X"00",X"A0",X"70",X"E8",X"B0",X"08",X"1F",X"00",X"3F",
		X"C0",X"2F",X"00",X"2F",X"40",X"0F",X"C0",X"0F",X"40",X"0F",X"00",X"3F",X"C0",X"0F",X"00",X"0F",
		X"40",X"1C",X"00",X"3C",X"C0",X"2C",X"00",X"2C",X"40",X"0C",X"C0",X"0C",X"40",X"0C",X"00",X"3C",
		X"C0",X"0C",X"00",X"0C",X"40",X"11",X"00",X"31",X"C0",X"21",X"00",X"21",X"40",X"01",X"C0",X"01",
		X"40",X"01",X"00",X"31",X"C0",X"01",X"00",X"01",X"40",X"CD",X"B0",X"3E",X"3A",X"00",X"50",X"CB",
		X"67",X"28",X"0A",X"21",X"AE",X"4C",X"CB",X"4E",X"20",X"03",X"3A",X"40",X"50",X"E6",X"0F",X"FE",
		X"0F",X"28",X"1B",X"0F",X"38",X"05",X"CD",X"4D",X"0F",X"18",X"13",X"0F",X"38",X"05",X"CD",X"99",
		X"0F",X"18",X"0B",X"0F",X"38",X"05",X"CD",X"80",X"0F",X"18",X"03",X"CD",X"35",X"0F",X"CD",X"C7",
		X"3C",X"CD",X"B2",X"0F",X"C9",X"3A",X"6A",X"4E",X"B7",X"C0",X"CD",X"6B",X"0F",X"B7",X"C8",X"3D",
		X"12",X"3C",X"CD",X"52",X"21",X"36",X"40",X"3E",X"10",X"32",X"6A",X"4E",X"C9",X"3A",X"6A",X"4E",
		X"B7",X"C0",X"CD",X"6B",X"0F",X"FE",X"02",X"28",X"0D",X"3C",X"12",X"CD",X"52",X"21",X"36",X"41",
		X"3E",X"10",X"32",X"6A",X"4E",X"C9",X"3D",X"32",X"AF",X"4C",X"C9",X"11",X"68",X"4E",X"1A",X"D6",
		X"05",X"ED",X"44",X"87",X"47",X"87",X"80",X"21",X"40",X"4E",X"CD",X"52",X"21",X"13",X"1A",X"C9",
		X"3A",X"6B",X"4E",X"B7",X"C0",X"CD",X"6B",X"0F",X"CD",X"52",X"21",X"7E",X"FE",X"5A",X"20",X"02",
		X"36",X"40",X"34",X"3E",X"10",X"32",X"6B",X"4E",X"C9",X"3A",X"6C",X"4E",X"B7",X"C0",X"CD",X"6B",
		X"0F",X"CD",X"52",X"21",X"7E",X"FE",X"41",X"20",X"02",X"36",X"5B",X"35",X"3E",X"10",X"32",X"6C",
		X"4E",X"C9",X"21",X"6A",X"4E",X"06",X"03",X"7E",X"B7",X"28",X"01",X"35",X"23",X"10",X"F8",X"C9",
		X"00",X"57",X"16",X"EB",X"21",X"3D",X"00",X"36",X"00",X"ED",X"53",X"43",X"02",X"ED",X"43",X"41",
		X"02",X"C1",X"E1",X"11",X"41",X"02",X"E5",X"C5",X"D5",X"0E",X"04",X"23",X"1A",X"BE",X"20",X"2C",
		X"13",X"0D",X"20",X"F7",X"78",X"D1",X"C1",X"D1",X"F6",X"80",X"E1",X"2B",X"2B",X"F5",X"7E",X"FE",
		X"27",X"28",X"01",X"23",X"F1",X"77",X"23",X"E5",X"2A",X"27",X"02",X"2B",X"7E",X"E1",X"22",X"65",
		X"21",X"6A",X"41",X"11",X"1D",X"00",X"3E",X"3F",X"0E",X"03",X"CD",X"A7",X"28",X"21",X"4A",X"42",
		X"0E",X"03",X"CD",X"A7",X"28",X"21",X"CA",X"41",X"06",X"03",X"36",X"3E",X"23",X"10",X"FB",X"21",
		X"2A",X"42",X"06",X"03",X"36",X"3D",X"23",X"10",X"FB",X"3E",X"1A",X"C3",X"30",X"10",X"3E",X"19",
		X"21",X"6A",X"45",X"11",X"1D",X"00",X"0E",X"04",X"CD",X"A7",X"28",X"21",X"2A",X"46",X"0E",X"04",
		X"C3",X"A7",X"28",X"21",X"83",X"4C",X"7E",X"B7",X"CA",X"29",X"10",X"FE",X"80",X"28",X"DF",X"C9",
		X"21",X"83",X"4C",X"34",X"C0",X"23",X"34",X"C9",X"E6",X"03",X"3C",X"47",X"0E",X"11",X"CB",X"09",
		X"10",X"FC",X"7E",X"B1",X"E6",X"0F",X"20",X"03",X"CB",X"01",X"C9",X"7E",X"B1",X"E6",X"0F",X"FE",
		X"09",X"C0",X"CB",X"01",X"C9",X"3A",X"83",X"4C",X"E6",X"0F",X"28",X"10",X"FE",X"03",X"C0",X"CD",
		X"D0",X"3A",X"C8",X"00",X"00",X"32",X"06",X"4E",X"32",X"20",X"4C",X"21",X"21",X"10",X"4E",X"11",
		X"08",X"4E",X"7E",X"B7",X"28",X"03",X"35",X"28",X"0D",X"EB",X"7E",X"B7",X"C8",X"35",X"C0",X"3A",
		X"06",X"4E",X"FE",X"03",X"D0",X"EB",X"AF",X"12",X"77",X"67",X"6F",X"22",X"EC",X"4F",X"22",X"CC",
		X"4F",X"3D",X"32",X"07",X"4E",X"CD",X"E0",X"31",X"3A",X"84",X"50",X"E6",X"C0",X"C9",X"3A",X"C6",
		X"50",X"E6",X"30",X"FE",X"30",X"C0",X"00",X"00",X"CD",X"6F",X"2E",X"35",X"21",X"03",X"4E",X"7E",
		X"FE",X"01",X"D8",X"21",X"07",X"4E",X"CB",X"46",X"C0",X"36",X"01",X"23",X"3E",X"FF",X"77",X"32",
		X"10",X"4E",X"CD",X"00",X"20",X"21",X"CC",X"4F",X"11",X"EC",X"4F",X"B7",X"28",X"0E",X"3D",X"28",
		X"17",X"3D",X"28",X"20",X"3D",X"28",X"3C",X"3D",X"28",X"45",X"18",X"4F",X"36",X"C0",X"23",X"36",
		X"07",X"EB",X"36",X"B8",X"23",X"36",X"50",X"C9",X"36",X"80",X"23",X"36",X"07",X"EB",X"36",X"48",
		X"23",X"36",X"48",X"C9",X"36",X"60",X"23",X"36",X"09",X"EB",X"36",X"C8",X"23",X"36",X"D8",X"3A",
		X"87",X"50",X"E6",X"C0",X"FE",X"C0",X"C9",X"3A",X"C9",X"50",X"E6",X"30",X"C8",X"FE",X"30",X"C8",
		X"00",X"00",X"E1",X"36",X"A0",X"23",X"36",X"07",X"EB",X"36",X"38",X"23",X"36",X"78",X"C9",X"36",
		X"40",X"23",X"36",X"16",X"EB",X"36",X"D8",X"23",X"36",X"28",X"C9",X"36",X"20",X"23",X"36",X"10",
		X"EB",X"36",X"48",X"23",X"36",X"A8",X"3A",X"8F",X"50",X"E6",X"C0",X"FE",X"40",X"C9",X"3A",X"C0",
		X"50",X"E6",X"30",X"C8",X"FE",X"20",X"C8",X"00",X"00",X"E5",X"3A",X"07",X"4E",X"E6",X"81",X"E8",
		X"CD",X"E3",X"11",X"21",X"E4",X"4F",X"11",X"EC",X"4F",X"CD",X"A2",X"2B",X"FE",X"04",X"D0",X"79",
		X"FE",X"04",X"D0",X"CD",X"00",X"20",X"01",X"09",X"CC",X"B7",X"28",X"1B",X"01",X"14",X"88",X"3D",
		X"28",X"15",X"01",X"09",X"68",X"3D",X"28",X"0F",X"01",X"07",X"A8",X"3D",X"28",X"09",X"01",X"09",
		X"CC",X"3D",X"28",X"03",X"01",X"19",X"24",X"21",X"CC",X"4F",X"70",X"23",X"71",X"21",X"07",X"4E",
		X"CB",X"FE",X"3E",X"1F",X"23",X"77",X"32",X"10",X"4E",X"21",X"00",X"01",X"11",X"02",X"4E",X"CD",
		X"29",X"3A",X"CD",X"39",X"3A",X"CD",X"F4",X"31",X"2A",X"C4",X"4F",X"E5",X"21",X"54",X"01",X"22",
		X"C4",X"4F",X"3A",X"83",X"4C",X"C6",X"60",X"47",X"3A",X"83",X"4C",X"B8",X"20",X"FA",X"E1",X"22",
		X"C4",X"4F",X"C9",X"3A",X"47",X"50",X"07",X"C9",X"3A",X"8E",X"50",X"E6",X"C0",X"C8",X"87",X"87",
		X"D8",X"00",X"00",X"C2",X"00",X"4E",X"3A",X"83",X"4C",X"E6",X"0F",X"C0",X"3A",X"07",X"4E",X"E6",
		X"03",X"E2",X"08",X"12",X"3E",X"FF",X"18",X"03",X"CD",X"00",X"20",X"21",X"83",X"4C",X"CB",X"66",
		X"28",X"3D",X"E6",X"87",X"F5",X"F5",X"CC",X"E5",X"28",X"F1",X"C4",X"B8",X"28",X"F1",X"3D",X"F5",
		X"F5",X"CC",X"34",X"29",X"F1",X"C4",X"10",X"29",X"F1",X"3D",X"F5",X"F5",X"CC",X"A8",X"29",X"F1",
		X"C4",X"62",X"29",X"F1",X"3D",X"F5",X"F5",X"CC",X"04",X"2A",X"F1",X"C4",X"B6",X"29",X"F1",X"3D",
		X"F5",X"F5",X"CC",X"66",X"2A",X"F1",X"C4",X"46",X"2A",X"F1",X"3D",X"C2",X"EC",X"22",X"C9",X"E6",
		X"87",X"F5",X"C4",X"DB",X"28",X"F1",X"3D",X"F5",X"C4",X"27",X"29",X"F1",X"3D",X"F5",X"C4",X"9F",
		X"29",X"F1",X"3D",X"F5",X"F5",X"CC",X"2A",X"2A",X"F1",X"C4",X"ED",X"29",X"F1",X"3D",X"F5",X"F5",
		X"CC",X"7D",X"2A",X"F1",X"C4",X"5D",X"2A",X"F1",X"3D",X"C2",X"EC",X"22",X"C9",X"3A",X"81",X"4C",
		X"FE",X"15",X"38",X"23",X"3A",X"83",X"4C",X"E6",X"3F",X"FE",X"13",X"20",X"1A",X"3A",X"D0",X"4C",
		X"21",X"DE",X"4C",X"BE",X"20",X"0D",X"23",X"34",X"C0",X"00",X"00",X"32",X"20",X"4C",X"3E",X"01",
		X"32",X"01",X"4C",X"77",X"23",X"36",X"00",X"21",X"03",X"4E",X"7E",X"FE",X"01",X"C0",X"23",X"7E",
		X"FE",X"34",X"D8",X"23",X"7E",X"FE",X"02",X"D8",X"3A",X"12",X"4E",X"B7",X"C0",X"CD",X"D7",X"3B",
		X"21",X"20",X"4C",X"CB",X"EE",X"C9",X"06",X"25",X"3E",X"82",X"32",X"5C",X"4C",X"C5",X"21",X"40",
		X"40",X"CD",X"DE",X"12",X"C1",X"10",X"F6",X"AF",X"3E",X"81",X"32",X"5C",X"4C",X"C9",X"E5",X"C5",
		X"ED",X"5F",X"CD",X"1F",X"13",X"8D",X"A0",X"20",X"21",X"7E",X"FE",X"FF",X"20",X"04",X"36",X"D7",
		X"18",X"13",X"FE",X"D4",X"20",X"09",X"E5",X"7C",X"C6",X"04",X"67",X"CD",X"40",X"1D",X"E1",X"CD",
		X"1F",X"13",X"20",X"06",X"35",X"3E",X"70",X"3D",X"20",X"FD",X"C1",X"7D",X"C6",X"20",X"6F",X"30",
		X"01",X"24",X"7C",X"FE",X"44",X"20",X"C8",X"E1",X"23",X"7D",X"FE",X"60",X"C8",X"18",X"BF",X"D6",
		X"D5",X"C8",X"3D",X"C8",X"3D",X"C8",X"C9",X"21",X"E4",X"4F",X"7E",X"E6",X"FE",X"57",X"23",X"7E",
		X"E6",X"FE",X"5F",X"2B",X"E5",X"CD",X"49",X"13",X"E1",X"78",X"B7",X"28",X"07",X"E5",X"7D",X"D6",
		X"30",X"6F",X"71",X"E1",X"CD",X"48",X"2D",X"18",X"E1",X"21",X"5F",X"13",X"06",X"14",X"7A",X"BE",
		X"23",X"20",X"07",X"7B",X"BE",X"23",X"20",X"03",X"4E",X"C9",X"23",X"23",X"10",X"F0",X"C9",X"70",
		X"98",X"00",X"70",X"C0",X"00",X"9C",X"98",X"00",X"9C",X"C0",X"00",X"88",X"4A",X"00",X"88",X"76",
		X"00",X"88",X"D8",X"00",X"88",X"7A",X"00",X"5A",X"60",X"00",X"B8",X"60",X"00",X"72",X"98",X"86",
		X"72",X"C0",X"86",X"9A",X"98",X"86",X"9A",X"C0",X"86",X"88",X"4C",X"89",X"88",X"74",X"89",X"88",
		X"D6",X"09",X"88",X"7C",X"09",X"5C",X"60",X"06",X"B6",X"60",X"06",X"DD",X"E5",X"E3",X"CD",X"AE",
		X"13",X"E3",X"DD",X"E1",X"C0",X"3A",X"B4",X"4F",X"87",X"D0",X"C8",X"33",X"33",X"C9",X"7C",X"FE",
		X"41",X"28",X"13",X"FE",X"42",X"C0",X"7D",X"D6",X"08",X"C8",X"3D",X"C8",X"D6",X"04",X"C8",X"3D",
		X"C8",X"D6",X"06",X"C8",X"3D",X"C9",X"7D",X"D6",X"E0",X"18",X"EC",X"4F",X"7D",X"D6",X"20",X"6F",
		X"7E",X"A6",X"79",X"C8",X"A6",X"C9",X"11",X"F2",X"4F",X"D9",X"11",X"62",X"50",X"06",X"02",X"CD",
		X"34",X"14",X"C4",X"5D",X"14",X"CD",X"3C",X"14",X"C4",X"5D",X"14",X"CD",X"44",X"14",X"C4",X"5D",
		X"14",X"21",X"E6",X"4F",X"CD",X"5D",X"14",X"CD",X"4C",X"14",X"CC",X"5D",X"14",X"21",X"E2",X"4F",
		X"CD",X"5D",X"14",X"CD",X"34",X"14",X"CC",X"5D",X"14",X"CD",X"3C",X"14",X"CC",X"5D",X"14",X"CD",
		X"44",X"14",X"CC",X"5D",X"14",X"CD",X"4C",X"14",X"C4",X"5D",X"14",X"3A",X"83",X"4C",X"47",X"E6",
		X"FC",X"FE",X"04",X"C0",X"78",X"2F",X"32",X"07",X"50",X"0F",X"D8",X"C3",X"B5",X"3A",X"B7",X"C8",
		X"2F",X"CB",X"7F",X"C9",X"3A",X"B4",X"4F",X"21",X"E4",X"4F",X"18",X"F2",X"3A",X"B8",X"4F",X"21",
		X"E8",X"4F",X"18",X"EA",X"3A",X"BA",X"4F",X"21",X"EA",X"4F",X"18",X"E2",X"21",X"EC",X"4F",X"3A",
		X"CC",X"4F",X"E6",X"FC",X"FE",X"AC",X"C8",X"FE",X"B0",X"C8",X"FE",X"B4",X"C9",X"E5",X"3A",X"20",
		X"4C",X"4F",X"3A",X"00",X"50",X"CB",X"67",X"20",X"02",X"CB",X"91",X"05",X"7E",X"23",X"CD",X"90",
		X"14",X"12",X"13",X"7E",X"CD",X"A3",X"14",X"12",X"13",X"E1",X"7D",X"D6",X"20",X"6F",X"7E",X"CB",
		X"51",X"28",X"02",X"EE",X"03",X"D9",X"12",X"13",X"D9",X"23",X"7E",X"D9",X"12",X"13",X"D9",X"C9",
		X"CB",X"51",X"20",X"07",X"CB",X"78",X"20",X"01",X"3D",X"3D",X"C9",X"2F",X"C6",X"10",X"CB",X"78",
		X"C0",X"3D",X"C9",X"CB",X"51",X"C8",X"2F",X"C6",X"11",X"C9",X"3A",X"B4",X"4F",X"07",X"30",X"09",
		X"21",X"E4",X"4F",X"CD",X"45",X"15",X"CD",X"14",X"15",X"3A",X"B8",X"4F",X"07",X"30",X"14",X"21",
		X"E8",X"4F",X"CD",X"45",X"15",X"3A",X"B4",X"4F",X"07",X"30",X"05",X"CD",X"21",X"15",X"18",X"03",
		X"CD",X"14",X"15",X"3A",X"BA",X"4F",X"07",X"D0",X"3A",X"B4",X"4F",X"07",X"30",X"0E",X"3A",X"B8",
		X"4F",X"07",X"38",X"1C",X"21",X"EA",X"4F",X"CD",X"45",X"15",X"18",X"35",X"3A",X"11",X"4E",X"B7",
		X"3A",X"B8",X"4F",X"28",X"13",X"07",X"38",X"08",X"21",X"EA",X"4F",X"CD",X"45",X"15",X"18",X"14",
		X"21",X"EA",X"4F",X"CD",X"45",X"15",X"18",X"2F",X"21",X"EA",X"4F",X"CD",X"45",X"15",X"3A",X"B8",
		X"4F",X"07",X"38",X"0D",X"ED",X"43",X"C2",X"4F",X"ED",X"53",X"E2",X"4F",X"01",X"00",X"00",X"50",
		X"58",X"3A",X"C6",X"4F",X"E6",X"F8",X"FE",X"B8",X"28",X"08",X"ED",X"43",X"C6",X"4F",X"ED",X"53",
		X"E6",X"4F",X"01",X"00",X"00",X"50",X"58",X"3A",X"10",X"4E",X"B7",X"C0",X"ED",X"43",X"CC",X"4F",
		X"ED",X"53",X"EC",X"4F",X"C9",X"11",X"00",X"00",X"42",X"4A",X"7E",X"FE",X"88",X"23",X"7E",X"20",
		X"12",X"FE",X"78",X"30",X"0E",X"FE",X"4A",X"38",X"0A",X"CD",X"7E",X"15",X"1E",X"88",X"3A",X"F5",
		X"45",X"47",X"C9",X"FE",X"98",X"20",X"0A",X"CD",X"9F",X"15",X"3A",X"EE",X"45",X"16",X"98",X"18",
		X"F0",X"FE",X"C0",X"C0",X"CD",X"9F",X"15",X"3A",X"E9",X"45",X"16",X"C0",X"18",X"E3",X"FE",X"72",
		X"30",X"41",X"FE",X"4E",X"38",X"3D",X"0E",X"B4",X"16",X"62",X"BA",X"D0",X"0E",X"94",X"15",X"BA",
		X"D0",X"0E",X"AC",X"15",X"BA",X"D0",X"0E",X"95",X"15",X"BA",X"D0",X"0E",X"B5",X"15",X"C9",X"2B",
		X"7E",X"FE",X"9A",X"30",X"1E",X"FE",X"76",X"38",X"1A",X"0E",X"B2",X"1E",X"8A",X"00",X"BB",X"D0",
		X"0E",X"92",X"1D",X"BB",X"D0",X"0E",X"AC",X"1D",X"BB",X"D0",X"0E",X"90",X"1D",X"BB",X"D0",X"0E",
		X"B0",X"1D",X"C9",X"33",X"33",X"C9",X"3A",X"01",X"4E",X"FE",X"10",X"3A",X"83",X"4C",X"E6",X"0F",
		X"FE",X"03",X"20",X"0A",X"CD",X"D0",X"3A",X"28",X"05",X"00",X"00",X"32",X"20",X"4C",X"21",X"E4",
		X"4F",X"7E",X"23",X"B6",X"E6",X"07",X"C0",X"2B",X"CD",X"7F",X"2C",X"7A",X"B7",X"28",X"06",X"FE",
		X"03",X"28",X"08",X"18",X"0A",X"7B",X"FE",X"40",X"D8",X"18",X"04",X"7B",X"FE",X"A0",X"D0",X"DD",
		X"21",X"00",X"40",X"DD",X"19",X"FD",X"21",X"00",X"44",X"FD",X"19",X"21",X"00",X"00",X"DD",X"56",
		X"E0",X"DD",X"5E",X"01",X"FD",X"46",X"E0",X"FD",X"4E",X"01",X"CD",X"88",X"16",X"DD",X"2B",X"FD",
		X"2B",X"DD",X"E5",X"E3",X"7D",X"FE",X"DF",X"20",X"0F",X"7C",X"FE",X"41",X"20",X"0A",X"11",X"20",
		X"00",X"19",X"FD",X"19",X"E3",X"CB",X"FD",X"E3",X"E3",X"DD",X"E1",X"DD",X"56",X"E0",X"DD",X"5E",
		X"FF",X"FD",X"46",X"E0",X"FD",X"4E",X"FF",X"CD",X"88",X"16",X"11",X"20",X"00",X"DD",X"19",X"FD",
		X"19",X"DD",X"56",X"FF",X"DD",X"5E",X"20",X"FD",X"46",X"FF",X"FD",X"4E",X"20",X"CD",X"88",X"16",
		X"DD",X"23",X"FD",X"23",X"CB",X"7D",X"28",X"09",X"CB",X"BD",X"11",X"E0",X"FF",X"DD",X"19",X"FD",
		X"19",X"DD",X"56",X"20",X"DD",X"5E",X"01",X"FD",X"46",X"20",X"FD",X"4E",X"01",X"CD",X"88",X"16",
		X"4D",X"55",X"21",X"05",X"4E",X"C3",X"C3",X"2A",X"24",X"CD",X"9B",X"13",X"7A",X"CD",X"B2",X"16",
		X"38",X"27",X"7B",X"CD",X"B2",X"16",X"38",X"21",X"7A",X"CD",X"DD",X"22",X"20",X"06",X"7B",X"CD",
		X"DD",X"22",X"28",X"43",X"78",X"CD",X"47",X"1D",X"28",X"0F",X"79",X"CD",X"47",X"1D",X"28",X"09",
		X"18",X"35",X"FE",X"D8",X"3F",X"D0",X"FE",X"E0",X"C9",X"DD",X"56",X"00",X"FD",X"46",X"00",X"CD",
		X"8A",X"21",X"7A",X"3C",X"20",X"07",X"78",X"CD",X"47",X"1D",X"C8",X"18",X"0A",X"7A",X"CD",X"DD",
		X"22",X"20",X"0D",X"DD",X"36",X"00",X"FF",X"78",X"CD",X"6D",X"1D",X"FD",X"77",X"00",X"2C",X"C9",
		X"78",X"CD",X"47",X"1D",X"C8",X"18",X"F0",X"DD",X"56",X"00",X"FD",X"46",X"00",X"CD",X"8A",X"21",
		X"78",X"CD",X"47",X"1D",X"C8",X"7A",X"3C",X"28",X"09",X"78",X"CD",X"6D",X"1D",X"FD",X"77",X"00",
		X"2C",X"C9",X"7C",X"CD",X"13",X"17",X"DD",X"70",X"00",X"FD",X"7E",X"00",X"CD",X"6D",X"1D",X"FD",
		X"77",X"00",X"C9",X"3D",X"06",X"CD",X"C8",X"05",X"3D",X"C8",X"06",X"CE",X"3D",X"C8",X"04",X"C9",
		X"21",X"20",X"4C",X"CB",X"EE",X"CD",X"C8",X"3F",X"C9",X"00",X"C4",X"AE",X"17",X"3A",X"3A",X"00",
		X"B7",X"28",X"07",X"CD",X"E4",X"11",X"AF",X"32",X"3A",X"00",X"36",X"08",X"CD",X"C1",X"17",X"CD",
		X"C1",X"17",X"21",X"95",X"02",X"CD",X"C4",X"17",X"3A",X"2A",X"00",X"DE",X"28",X"DE",X"08",X"38",
		X"03",X"CD",X"BE",X"13",X"21",X"C1",X"02",X"CD",X"C4",X"17",X"21",X"82",X"01",X"34",X"7E",X"CD",
		X"98",X"17",X"CD",X"C1",X"17",X"3A",X"89",X"02",X"B7",X"28",X"14",X"21",X"12",X"00",X"22",X"54",
		X"00",X"21",X"29",X"02",X"D5",X"CD",X"5C",X"0A",X"D1",X"21",X"94",X"17",X"CD",X"C4",X"17",X"21",
		X"83",X"01",X"CD",X"BE",X"17",X"21",X"D4",X"01",X"CD",X"BE",X"17",X"CD",X"C1",X"17",X"CD",X"C1",
		X"17",X"C3",X"12",X"17",X"03",X"20",X"2D",X"20",X"D5",X"C5",X"16",X"00",X"06",X"64",X"CD",X"D1",
		X"17",X"06",X"0A",X"CD",X"D1",X"17",X"06",X"01",X"CD",X"D1",X"17",X"C1",X"D1",X"C9",X"E5",X"21",
		X"46",X"00",X"3A",X"47",X"00",X"3D",X"BE",X"D4",X"08",X"17",X"30",X"FA",X"E1",X"C9",X"CD",X"C4",
		X"17",X"21",X"C7",X"02",X"7E",X"B7",X"C8",X"23",X"4E",X"F5",X"CD",X"12",X"00",X"F1",X"3D",X"18",
		X"F5",X"0E",X"30",X"90",X"38",X"03",X"0C",X"18",X"FA",X"80",X"F5",X"79",X"FE",X"30",X"20",X"04",
		X"7A",X"B7",X"28",X"05",X"CD",X"12",X"00",X"16",X"01",X"F1",X"C9",X"AF",X"00",X"00",X"3E",X"01",
		X"18",X"02",X"3E",X"02",X"C5",X"D5",X"C5",X"4F",X"ED",X"5B",X"2D",X"02",X"2A",X"27",X"02",X"B9",
		X"3E",X"01",X"32",X"04",X"50",X"21",X"D0",X"4C",X"34",X"7E",X"FE",X"3C",X"D8",X"36",X"00",X"23",
		X"34",X"7E",X"FE",X"1E",X"D8",X"AF",X"77",X"32",X"04",X"50",X"C9",X"3A",X"83",X"4C",X"FE",X"01",
		X"20",X"0A",X"CC",X"D0",X"3A",X"28",X"05",X"00",X"00",X"32",X"20",X"4C",X"CD",X"DD",X"18",X"CD",
		X"8E",X"18",X"D5",X"3A",X"03",X"4E",X"3D",X"28",X"0E",X"3A",X"06",X"4E",X"FE",X"01",X"30",X"07",
		X"3A",X"04",X"4E",X"FE",X"10",X"38",X"11",X"CD",X"B4",X"1A",X"20",X"0C",X"7E",X"CD",X"FE",X"18",
		X"28",X"06",X"CD",X"D3",X"18",X"CD",X"07",X"19",X"E1",X"3A",X"03",X"4E",X"3D",X"28",X"10",X"3A",
		X"06",X"4E",X"FE",X"01",X"06",X"20",X"38",X"02",X"06",X"10",X"3A",X"04",X"4E",X"B8",X"D8",X"CD",
		X"B4",X"1A",X"C0",X"7E",X"CD",X"FE",X"18",X"C8",X"CD",X"D3",X"18",X"E5",X"CD",X"5C",X"19",X"E1",
		X"20",X"09",X"E5",X"CD",X"61",X"19",X"E1",X"C8",X"79",X"D7",X"4F",X"C3",X"07",X"19",X"11",X"E4",
		X"4F",X"21",X"E8",X"4F",X"CD",X"42",X"19",X"13",X"23",X"47",X"CD",X"42",X"19",X"80",X"47",X"2E",
		X"EB",X"CD",X"42",X"19",X"2B",X"1B",X"4F",X"CD",X"42",X"19",X"81",X"1E",X"DA",X"2E",X"D8",X"B8",
		X"D0",X"EB",X"3A",X"00",X"50",X"0F",X"D8",X"3A",X"55",X"50",X"07",X"C9",X"3A",X"87",X"50",X"E6",
		X"C0",X"C8",X"07",X"07",X"D8",X"00",X"00",X"21",X"12",X"4E",X"3A",X"40",X"50",X"34",X"D8",X"21",
		X"03",X"4E",X"35",X"E5",X"7D",X"C6",X"10",X"6F",X"CD",X"1C",X"19",X"E1",X"C9",X"21",X"EC",X"4F",
		X"3A",X"DC",X"4F",X"CD",X"FE",X"18",X"C8",X"CD",X"14",X"1C",X"30",X"05",X"CD",X"34",X"1C",X"18",
		X"08",X"E5",X"CD",X"6F",X"19",X"E1",X"CD",X"1F",X"19",X"2E",X"DC",X"C3",X"07",X"19",X"D7",X"E6",
		X"0F",X"FE",X"06",X"C8",X"FE",X"09",X"C9",X"7E",X"D7",X"E6",X"0F",X"E5",X"CD",X"F6",X"19",X"E1",
		X"47",X"79",X"A0",X"20",X"04",X"79",X"D7",X"A0",X"C8",X"23",X"77",X"C9",X"11",X"E4",X"4F",X"CD",
		X"42",X"19",X"47",X"23",X"13",X"CD",X"42",X"19",X"B8",X"30",X"0B",X"CD",X"48",X"19",X"D7",X"47",
		X"CD",X"51",X"19",X"B0",X"4F",X"C9",X"CD",X"51",X"19",X"D7",X"47",X"23",X"13",X"CD",X"48",X"19",
		X"18",X"F1",X"1A",X"96",X"F0",X"ED",X"44",X"C9",X"1A",X"96",X"C8",X"3E",X"08",X"D8",X"3E",X"01",
		X"C9",X"2B",X"1B",X"1A",X"96",X"C8",X"3E",X"04",X"D8",X"3E",X"02",X"C9",X"11",X"E8",X"4F",X"18",
		X"03",X"11",X"E4",X"4F",X"21",X"EA",X"4F",X"1A",X"BE",X"C8",X"23",X"13",X"1A",X"BE",X"C9",X"CD",
		X"94",X"19",X"D8",X"3A",X"8E",X"50",X"E6",X"C0",X"18",X"12",X"3A",X"FF",X"50",X"E6",X"30",X"FE",
		X"30",X"20",X"09",X"00",X"00",X"ED",X"5B",X"EC",X"4F",X"32",X"03",X"4E",X"ED",X"53",X"E0",X"4F",
		X"11",X"E0",X"4F",X"C9",X"11",X"E8",X"4F",X"3A",X"07",X"4E",X"E6",X"81",X"37",X"E8",X"3A",X"10",
		X"4E",X"07",X"D8",X"07",X"D8",X"CD",X"00",X"20",X"87",X"21",X"B4",X"19",X"CD",X"52",X"21",X"5E",
		X"23",X"56",X"AF",X"C9",X"C8",X"50",X"58",X"50",X"B8",X"D8",X"48",X"78",X"C8",X"20",X"58",X"B0",
		X"3A",X"07",X"4E",X"E6",X"81",X"E8",X"3A",X"10",X"4E",X"07",X"D8",X"07",X"D8",X"CD",X"00",X"20",
		X"87",X"21",X"B4",X"19",X"CD",X"52",X"21",X"11",X"EC",X"4F",X"1A",X"BE",X"C0",X"23",X"13",X"1A",
		X"BE",X"C0",X"AF",X"32",X"08",X"4E",X"32",X"10",X"4E",X"67",X"6F",X"22",X"EC",X"4F",X"22",X"CC",
		X"4F",X"3D",X"32",X"07",X"4E",X"C9",X"F5",X"7D",X"C6",X"10",X"6F",X"56",X"23",X"5E",X"3A",X"E4",
		X"4F",X"FE",X"88",X"21",X"5A",X"1A",X"06",X"0B",X"28",X"20",X"3A",X"E5",X"4F",X"FE",X"C0",X"21",
		X"8D",X"1A",X"06",X"0A",X"28",X"29",X"21",X"99",X"1A",X"06",X"09",X"FE",X"98",X"28",X"20",X"21",
		X"6F",X"1A",X"06",X"08",X"FE",X"60",X"28",X"0F",X"F1",X"C9",X"3A",X"11",X"4E",X"B7",X"28",X"0F",
		X"21",X"54",X"1A",X"06",X"0D",X"18",X"08",X"3A",X"11",X"4E",X"B7",X"28",X"02",X"06",X"0A",X"7A",
		X"BE",X"23",X"20",X"06",X"7B",X"BE",X"23",X"28",X"07",X"2B",X"23",X"23",X"10",X"F1",X"F1",X"C9",
		X"46",X"F1",X"A0",X"C9",X"88",X"78",X"0E",X"88",X"D8",X"07",X"58",X"D8",X"07",X"B8",X"D8",X"07",
		X"68",X"78",X"0E",X"B8",X"78",X"0E",X"48",X"60",X"0D",X"58",X"60",X"0D",X"B8",X"60",X"0B",X"58",
		X"C0",X"0D",X"B8",X"C0",X"0B",X"68",X"98",X"0D",X"B8",X"98",X"0B",X"48",X"78",X"0D",X"88",X"78",
		X"07",X"B8",X"78",X"0B",X"88",X"38",X"0E",X"58",X"60",X"0D",X"B8",X"98",X"0B",X"88",X"D8",X"07",
		X"58",X"98",X"0D",X"68",X"98",X"0D",X"B8",X"98",X"0B",X"68",X"78",X"0D",X"88",X"78",X"0E",X"B8",
		X"78",X"0B",X"48",X"60",X"0D",X"58",X"60",X"0D",X"B8",X"60",X"0B",X"88",X"D8",X"07",X"58",X"C0",
		X"0D",X"B0",X"C0",X"0B",X"E5",X"7D",X"C6",X"10",X"6F",X"CD",X"BE",X"1A",X"E1",X"C9",X"7E",X"23",
		X"B6",X"2B",X"E6",X"07",X"C9",X"3A",X"06",X"4E",X"FE",X"01",X"30",X"06",X"3A",X"0F",X"4E",X"FE",
		X"01",X"D8",X"79",X"E6",X"06",X"79",X"28",X"04",X"EE",X"06",X"4F",X"C9",X"EE",X"09",X"4F",X"C9",
		X"3A",X"20",X"4C",X"CB",X"57",X"28",X"1F",X"3A",X"83",X"4C",X"E6",X"3F",X"FE",X"31",X"20",X"16",
		X"3A",X"D0",X"4C",X"21",X"DA",X"4C",X"BE",X"20",X"09",X"23",X"34",X"20",X"09",X"00",X"00",X"22",
		X"1F",X"4C",X"77",X"23",X"36",X"00",X"11",X"E4",X"4F",X"21",X"E8",X"4F",X"D5",X"CD",X"14",X"1B",
		X"D1",X"21",X"EA",X"4F",X"E5",X"CD",X"33",X"1B",X"E1",X"79",X"B7",X"C8",X"7D",X"D6",X"10",X"6F",
		X"7E",X"CD",X"FE",X"18",X"C8",X"7E",X"D7",X"E6",X"0F",X"57",X"A1",X"20",X"03",X"7A",X"A0",X"C8",
		X"23",X"77",X"C9",X"01",X"00",X"00",X"CD",X"BE",X"1A",X"C0",X"1A",X"FE",X"50",X"38",X"1B",X"FE",
		X"C0",X"30",X"31",X"13",X"1A",X"FE",X"40",X"38",X"0A",X"FE",X"D0",X"D8",X"23",X"7E",X"FE",X"40",
		X"D0",X"18",X"4B",X"23",X"7E",X"FE",X"D0",X"D8",X"18",X"44",X"7E",X"FE",X"C0",X"D8",X"23",X"13",
		X"1A",X"FE",X"90",X"7E",X"38",X"07",X"FE",X"B0",X"D8",X"16",X"C0",X"18",X"21",X"FE",X"B0",X"D0",
		X"16",X"60",X"18",X"1A",X"7E",X"FE",X"50",X"D0",X"23",X"13",X"1A",X"FE",X"B0",X"7E",X"38",X"07",
		X"FE",X"90",X"D8",X"16",X"C0",X"18",X"07",X"FE",X"90",X"D0",X"16",X"60",X"18",X"00",X"7E",X"BA",
		X"0E",X"01",X"D8",X"06",X"08",X"2B",X"7E",X"07",X"0E",X"02",X"D8",X"0E",X"04",X"C9",X"2B",X"7E",
		X"FE",X"88",X"0E",X"02",X"D8",X"06",X"04",X"23",X"7E",X"07",X"0E",X"01",X"D8",X"0E",X"08",X"C9",
		X"21",X"E8",X"4F",X"11",X"F0",X"4F",X"1A",X"3C",X"28",X"0A",X"12",X"36",X"A0",X"D5",X"E5",X"CD",
		X"CD",X"1B",X"E1",X"D1",X"13",X"1A",X"3C",X"C8",X"12",X"23",X"23",X"36",X"70",X"23",X"36",X"B0",
		X"1A",X"3C",X"C0",X"7D",X"D6",X"21",X"6F",X"36",X"E0",X"23",X"36",X"07",X"7D",X"FE",X"C9",X"CA",
		X"6C",X"39",X"36",X"05",X"C3",X"79",X"39",X"3A",X"80",X"50",X"F5",X"0F",X"0F",X"E6",X"03",X"06",
		X"03",X"28",X"09",X"04",X"3D",X"28",X"05",X"04",X"3D",X"28",X"01",X"04",X"78",X"32",X"01",X"4C",
		X"F1",X"E6",X"C0",X"FE",X"40",X"C9",X"3A",X"CC",X"50",X"E6",X"30",X"C8",X"FE",X"20",X"C8",X"00",
		X"00",X"32",X"19",X"4E",X"11",X"E4",X"4F",X"3A",X"06",X"4E",X"FE",X"01",X"3F",X"D0",X"1A",X"96",
		X"30",X"02",X"ED",X"44",X"FE",X"48",X"D0",X"23",X"13",X"1A",X"96",X"2B",X"1B",X"30",X"02",X"ED",
		X"44",X"FE",X"48",X"C9",X"1A",X"96",X"0E",X"24",X"C8",X"23",X"13",X"1A",X"96",X"0E",X"18",X"C8",
		X"2B",X"1B",X"CD",X"1C",X"19",X"79",X"06",X"09",X"A0",X"20",X"02",X"06",X"06",X"79",X"A8",X"4F",
		X"06",X"90",X"A0",X"20",X"02",X"06",X"60",X"79",X"A8",X"4F",X"C9",X"21",X"E8",X"4F",X"CD",X"64",
		X"1C",X"21",X"EA",X"4F",X"11",X"E4",X"4F",X"1A",X"13",X"FE",X"58",X"28",X"1A",X"FE",X"C8",X"C0",
		X"1A",X"FE",X"61",X"D0",X"7E",X"FE",X"B8",X"C0",X"23",X"7E",X"FE",X"C0",X"28",X"1A",X"FE",X"98",
		X"28",X"16",X"FE",X"78",X"C0",X"18",X"11",X"1A",X"FE",X"61",X"D0",X"7E",X"FE",X"48",X"C0",X"23",
		X"7E",X"FE",X"78",X"28",X"03",X"FE",X"98",X"C0",X"7D",X"D6",X"10",X"6F",X"36",X"08",X"C9",X"3A",
		X"C0",X"50",X"E6",X"1F",X"FE",X"1F",X"0E",X"FF",X"C9",X"06",X"3A",X"80",X"50",X"E6",X"C0",X"C8",
		X"F3",X"CD",X"66",X"0B",X"18",X"FB",X"CD",X"8C",X"1D",X"FE",X"06",X"38",X"02",X"3E",X"05",X"87",
		X"87",X"21",X"11",X"1D",X"CD",X"52",X"21",X"7E",X"4F",X"E5",X"C5",X"CD",X"29",X"1D",X"C1",X"E1",
		X"79",X"20",X"05",X"CC",X"77",X"1D",X"18",X"0D",X"3A",X"06",X"4E",X"FE",X"05",X"38",X"05",X"E6",
		X"03",X"28",X"01",X"0D",X"79",X"32",X"CE",X"4F",X"23",X"7E",X"32",X"92",X"4C",X"23",X"7E",X"32",
		X"94",X"4C",X"23",X"7E",X"32",X"96",X"4C",X"3A",X"81",X"4C",X"FE",X"10",X"D8",X"3A",X"83",X"4C",
		X"FE",X"09",X"C0",X"CD",X"D0",X"3A",X"C8",X"00",X"00",X"32",X"19",X"4E",X"AF",X"32",X"03",X"4E",
		X"C9",X"0F",X"0E",X"0E",X"0C",X"80",X"0F",X"0F",X"0D",X"82",X"81",X"81",X"0F",X"84",X"83",X"83",
		X"81",X"86",X"85",X"85",X"83",X"89",X"88",X"88",X"85",X"21",X"E4",X"4F",X"CD",X"7F",X"2C",X"21",
		X"00",X"40",X"19",X"7E",X"2B",X"A6",X"F5",X"CD",X"50",X"21",X"F1",X"A6",X"23",X"A6",X"3C",X"C9",
		X"7E",X"E6",X"E0",X"F6",X"03",X"77",X"C9",X"E6",X"1F",X"FE",X"06",X"C8",X"FE",X"02",X"C8",X"FE",
		X"04",X"C9",X"3A",X"06",X"4E",X"FE",X"03",X"38",X"04",X"D6",X"03",X"18",X"F8",X"3C",X"FE",X"03",
		X"20",X"01",X"3C",X"32",X"19",X"4E",X"FE",X"01",X"C0",X"3E",X"06",X"18",X"F6",X"E6",X"E0",X"C5",
		X"47",X"3A",X"19",X"4E",X"B0",X"C1",X"C9",X"3D",X"F5",X"3A",X"80",X"50",X"CB",X"67",X"18",X"07",
		X"3A",X"06",X"4E",X"FE",X"01",X"38",X"03",X"F1",X"3D",X"C9",X"F1",X"C9",X"3A",X"06",X"4E",X"FE",
		X"05",X"D0",X"FE",X"02",X"D8",X"F5",X"3A",X"03",X"4E",X"B7",X"28",X"0A",X"3A",X"04",X"4E",X"FE",
		X"10",X"38",X"03",X"F1",X"3C",X"C9",X"F1",X"C9",X"21",X"40",X"4E",X"0E",X"05",X"06",X"03",X"36",
		X"4B",X"23",X"36",X"52",X"23",X"36",X"4C",X"23",X"23",X"23",X"23",X"0D",X"20",X"EF",X"3E",X"81",
		X"32",X"AC",X"4C",X"C9",X"21",X"AE",X"4C",X"7E",X"B7",X"C8",X"CB",X"57",X"28",X"0B",X"CB",X"96",
		X"E5",X"CD",X"F1",X"1D",X"E1",X"ED",X"43",X"66",X"4E",X"ED",X"4B",X"66",X"4E",X"78",X"B1",X"20",
		X"03",X"36",X"00",X"C9",X"7E",X"E6",X"82",X"C2",X"52",X"3D",X"7E",X"E6",X"41",X"C2",X"6F",X"3D",
		X"C9",X"11",X"00",X"4D",X"21",X"80",X"4D",X"01",X"00",X"00",X"CD",X"64",X"1E",X"38",X"09",X"CD",
		X"1D",X"1E",X"78",X"B7",X"C8",X"C3",X"11",X"1E",X"CD",X"11",X"1E",X"79",X"B7",X"C8",X"C3",X"1D",
		X"1E",X"11",X"80",X"4D",X"C5",X"41",X"CD",X"20",X"1E",X"78",X"C1",X"4F",X"C9",X"11",X"00",X"4D",
		X"21",X"5E",X"4E",X"C5",X"06",X"03",X"36",X"40",X"23",X"10",X"FB",X"06",X"03",X"1A",X"77",X"23",
		X"13",X"10",X"FA",X"C1",X"21",X"5B",X"4E",X"11",X"61",X"4E",X"CD",X"64",X"1E",X"D8",X"C8",X"7D",
		X"D6",X"03",X"6F",X"7B",X"D6",X"03",X"5F",X"C5",X"06",X"06",X"1A",X"F5",X"7E",X"12",X"F1",X"77",
		X"23",X"13",X"10",X"F6",X"C1",X"04",X"78",X"FE",X"05",X"C8",X"7B",X"D6",X"09",X"5F",X"7D",X"D6",
		X"09",X"6F",X"18",X"D6",X"E5",X"D5",X"CD",X"6C",X"1E",X"D1",X"E1",X"C9",X"1A",X"BE",X"D8",X"C0",
		X"13",X"23",X"1A",X"BE",X"D8",X"C0",X"13",X"23",X"1A",X"BE",X"C9",X"00",X"23",X"F6",X"01",X"C9",
		X"E3",X"E1",X"D5",X"7E",X"23",X"E6",X"03",X"FE",X"02",X"20",X"06",X"5E",X"23",X"56",X"2B",X"18",
		X"03",X"11",X"03",X"00",X"19",X"D1",X"18",X"B3",X"21",X"10",X"00",X"E5",X"3A",X"29",X"00",X"32",
		X"40",X"02",X"AF",X"32",X"28",X"00",X"CD",X"AF",X"14",X"DA",X"BD",X"1F",X"CD",X"EC",X"16",X"38",
		X"77",X"CD",X"57",X"16",X"CD",X"AF",X"14",X"FE",X"23",X"20",X"06",X"CD",X"CA",X"13",X"CD",X"E4",
		X"15",X"D5",X"3A",X"2F",X"02",X"B7",X"20",X"07",X"CD",X"22",X"15",X"38",X"31",X"18",X"0C",X"CD",
		X"26",X"15",X"30",X"4D",X"2A",X"40",X"00",X"7C",X"B5",X"28",X"23",X"CB",X"66",X"28",X"3A",X"CB",
		X"5E",X"C4",X"25",X"1B",X"CD",X"59",X"18",X"D1",X"CA",X"C5",X"1F",X"3A",X"28",X"00",X"B7",X"28",
		X"04",X"B9",X"C4",X"0D",X"1B",X"79",X"32",X"28",X"00",X"0E",X"01",X"C3",X"C5",X"1F",X"2A",X"3E",
		X"00",X"7C",X"B5",X"28",X"0D",X"23",X"23",X"5E",X"23",X"56",X"EB",X"AF",X"47",X"4F",X"D1",X"C3",
		X"C5",X"1F",X"3A",X"81",X"00",X"3D",X"C4",X"EE",X"17",X"CD",X"19",X"1B",X"21",X"00",X"00",X"18",
		X"EA",X"D1",X"CD",X"20",X"19",X"C3",X"A6",X"1E",X"21",X"40",X"02",X"FE",X"30",X"38",X"0B",X"FE",
		X"3A",X"30",X"07",X"7E",X"CD",X"96",X"21",X"C3",X"C5",X"1F",X"1A",X"FE",X"22",X"28",X"04",X"FE",
		X"27",X"20",X"21",X"47",X"21",X"00",X"00",X"E5",X"CD",X"CA",X"13",X"B8",X"20",X"06",X"CD",X"CA",
		X"13",X"B8",X"20",X"0D",X"FE",X"0D",X"20",X"05",X"CD",X"15",X"1B",X"18",X"04",X"65",X"6F",X"18",
		X"E7",X"C1",X"18",X"61",X"FE",X"5E",X"20",X"20",X"7E",X"3D",X"07",X"07",X"07",X"07",X"F6",X"17",
		X"4F",X"06",X"0F",X"C5",X"CD",X"CA",X"13",X"CD",X"FF",X"16",X"E5",X"21",X"2C",X"22",X"CD",X"59",
		X"21",X"38",X"2C",X"7E",X"E1",X"77",X"18",X"73",X"FE",X"2B",X"28",X"6F",X"FE",X"28",X"20",X"0D",
		X"3A",X"28",X"00",X"F5",X"AF",X"32",X"28",X"00",X"01",X"11",X"0D",X"18",X"5D",X"FE",X"2D",X"20",
		X"05",X"01",X"18",X"0E",X"18",X"54",X"FE",X"23",X"20",X"06",X"01",X"15",X"0C",X"18",X"4B",X"E1",
		X"CD",X"01",X"1B",X"18",X"46",X"CD",X"01",X"1B",X"01",X"00",X"00",X"18",X"2D",X"CD",X"01",X"1B",
		X"01",X"00",X"00",X"60",X"68",X"22",X"3C",X"02",X"ED",X"43",X"3E",X"02",X"CD",X"AF",X"14",X"21",
		X"39",X"22",X"CD",X"59",X"21",X"30",X"12",X"CD",X"EC",X"16",X"38",X"D9",X"CD",X"57",X"16",X"CD",
		X"26",X"15",X"38",X"D1",X"CD",X"20",X"19",X"18",X"E3",X"4E",X"E1",X"7D",X"E6",X"0F",X"B9",X"30",
		X"10",X"E5",X"2A",X"3C",X"02",X"E5",X"2A",X"3E",X"02",X"E5",X"C5",X"CD",X"CA",X"13",X"C3",X"32",
		X"3A",X"06",X"4E",X"FE",X"06",X"D8",X"D6",X"06",X"18",X"F9",X"3A",X"07",X"4E",X"E6",X"81",X"E8",
		X"CD",X"D7",X"31",X"3A",X"12",X"4E",X"FE",X"55",X"38",X"17",X"3A",X"20",X"4C",X"CB",X"57",X"C0",
		X"3A",X"83",X"4C",X"E6",X"FD",X"FE",X"05",X"C0",X"CD",X"D0",X"3A",X"C8",X"00",X"00",X"32",X"12",
		X"4E",X"21",X"EC",X"4F",X"7E",X"23",X"B6",X"2B",X"E6",X"07",X"C0",X"CD",X"00",X"20",X"5F",X"FE",
		X"03",X"28",X"06",X"D5",X"CD",X"57",X"21",X"D1",X"D8",X"3A",X"DC",X"4F",X"CD",X"C0",X"20",X"7B",
		X"87",X"87",X"81",X"87",X"21",X"6D",X"20",X"CD",X"64",X"20",X"CD",X"9D",X"20",X"21",X"12",X"4E",
		X"7E",X"82",X"77",X"C9",X"85",X"6F",X"30",X"01",X"24",X"46",X"23",X"4E",X"C9",X"A7",X"A7",X"A7",
		X"A7",X"A7",X"A7",X"A7",X"A7",X"A9",X"A9",X"A8",X"A8",X"A8",X"A8",X"A9",X"A9",X"AA",X"AB",X"AA",
		X"AB",X"AA",X"AB",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"AE",X"AF",X"AC",X"AD",X"B8",X"B9",X"B8",
		X"B9",X"B8",X"B9",X"B8",X"B9",X"B2",X"B3",X"B5",X"B4",X"B0",X"B1",X"B7",X"B6",X"21",X"EC",X"4F",
		X"D5",X"C5",X"CD",X"7F",X"2C",X"21",X"00",X"40",X"19",X"C1",X"D1",X"16",X"00",X"7B",X"FE",X"03",
		X"28",X"26",X"CD",X"CA",X"20",X"7D",X"C6",X"1F",X"6F",X"30",X"01",X"24",X"41",X"C3",X"CA",X"20",
		X"0E",X"00",X"E6",X"0F",X"C8",X"0F",X"D8",X"0C",X"18",X"FB",X"7E",X"FE",X"FF",X"20",X"03",X"70",
		X"14",X"C9",X"CD",X"74",X"21",X"D0",X"70",X"C9",X"3A",X"DC",X"4F",X"0F",X"38",X"41",X"0F",X"38",
		X"2D",X"0F",X"38",X"16",X"0F",X"D0",X"2B",X"3E",X"AE",X"01",X"AC",X"BB",X"CD",X"32",X"21",X"CD",
		X"50",X"21",X"3E",X"AE",X"01",X"AD",X"BD",X"C3",X"32",X"21",X"CD",X"50",X"21",X"3E",X"AC",X"01",
		X"AE",X"BB",X"CD",X"32",X"21",X"2B",X"3E",X"AC",X"01",X"AF",X"BA",X"C3",X"32",X"21",X"3E",X"AD",
		X"01",X"AE",X"BD",X"CD",X"32",X"21",X"2B",X"3E",X"AD",X"01",X"AF",X"BC",X"C3",X"32",X"21",X"3E",
		X"AF",X"01",X"AC",X"BA",X"CD",X"32",X"21",X"CD",X"50",X"21",X"3E",X"AF",X"01",X"AD",X"BC",X"C3",
		X"32",X"21",X"BE",X"20",X"02",X"70",X"C9",X"3E",X"FF",X"BE",X"C0",X"71",X"14",X"3A",X"77",X"50",
		X"87",X"C9",X"10",X"03",X"00",X"E6",X"C0",X"C8",X"87",X"87",X"D8",X"00",X"00",X"14",X"77",X"C9",
		X"3E",X"20",X"85",X"6F",X"D0",X"24",X"C9",X"CD",X"7F",X"2C",X"21",X"00",X"40",X"19",X"CD",X"74",
		X"21",X"D8",X"2B",X"CD",X"74",X"21",X"D8",X"11",X"20",X"00",X"19",X"CD",X"74",X"21",X"D8",X"23",
		X"CD",X"74",X"21",X"C9",X"7E",X"FE",X"BE",X"D0",X"FE",X"A7",X"3F",X"C9",X"7A",X"FE",X"BE",X"30",
		X"06",X"FE",X"A7",X"38",X"02",X"AF",X"C9",X"F6",X"FF",X"C9",X"7A",X"CD",X"75",X"21",X"D0",X"3A",
		X"12",X"4E",X"3D",X"32",X"12",X"4E",X"16",X"FF",X"DD",X"72",X"00",X"E5",X"D5",X"21",X"01",X"00",
		X"11",X"02",X"4E",X"CD",X"29",X"3A",X"CD",X"C0",X"31",X"D1",X"E1",X"C9",X"3A",X"81",X"4C",X"FE",
		X"20",X"38",X"1F",X"3A",X"83",X"4C",X"E6",X"3F",X"FE",X"35",X"20",X"16",X"3A",X"D0",X"4C",X"21",
		X"D8",X"4C",X"BE",X"20",X"08",X"23",X"34",X"C0",X"00",X"00",X"32",X"20",X"4C",X"77",X"23",X"36",
		X"00",X"00",X"21",X"12",X"40",X"06",X"0C",X"CD",X"66",X"23",X"21",X"5F",X"42",X"11",X"20",X"00",
		X"06",X"07",X"36",X"F7",X"19",X"10",X"FB",X"06",X"05",X"36",X"40",X"19",X"10",X"FB",X"21",X"1D",
		X"40",X"11",X"BF",X"43",X"01",X"E0",X"FF",X"3A",X"20",X"4C",X"CB",X"57",X"3A",X"1C",X"4C",X"28",
		X"03",X"3A",X"1D",X"4C",X"3D",X"F8",X"C8",X"FE",X"06",X"38",X"02",X"3E",X"06",X"F5",X"36",X"C8",
		X"2B",X"36",X"C9",X"2B",X"EB",X"36",X"CA",X"09",X"36",X"CB",X"09",X"EB",X"3D",X"20",X"EF",X"21",
		X"BF",X"47",X"11",X"1D",X"44",X"F1",X"08",X"3E",X"01",X"77",X"09",X"77",X"09",X"EB",X"77",X"2B",
		X"77",X"2B",X"EB",X"08",X"3D",X"C8",X"18",X"EE",X"CD",X"44",X"23",X"3A",X"9F",X"4C",X"B7",X"C8",
		X"FE",X"06",X"38",X"02",X"3E",X"06",X"01",X"20",X"00",X"21",X"5F",X"40",X"D9",X"21",X"22",X"40",
		X"11",X"02",X"40",X"36",X"C2",X"23",X"36",X"C3",X"23",X"EB",X"36",X"C4",X"23",X"36",X"C5",X"23",
		X"EB",X"D9",X"36",X"C6",X"09",X"36",X"C7",X"09",X"D9",X"3D",X"20",X"E7",X"01",X"9C",X"22",X"3A",
		X"9F",X"4C",X"F5",X"FE",X"13",X"38",X"02",X"3E",X"13",X"81",X"4F",X"30",X"01",X"04",X"F1",X"FE",
		X"06",X"38",X"02",X"3E",X"06",X"21",X"22",X"44",X"11",X"02",X"44",X"08",X"0A",X"77",X"23",X"77",
		X"23",X"EB",X"77",X"23",X"77",X"23",X"EB",X"03",X"08",X"3D",X"20",X"EF",X"C9",X"07",X"07",X"07",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"0F",X"0F",X"11",X"11",X"12",X"12",X"14",X"14",X"05",
		X"05",X"05",X"05",X"05",X"05",X"CD",X"CF",X"22",X"C4",X"7C",X"21",X"C4",X"0D",X"3C",X"C0",X"53",
		X"CD",X"CF",X"22",X"C4",X"7C",X"21",X"C4",X"0D",X"3C",X"C0",X"CB",X"E1",X"33",X"33",X"C9",X"7A",
		X"D6",X"FC",X"C8",X"3D",X"C8",X"3D",X"C8",X"3D",X"C8",X"7A",X"FE",X"D2",X"C8",X"D6",X"CC",X"C8",
		X"3D",X"C8",X"3D",X"C8",X"3D",X"C9",X"BA",X"C0",X"BB",X"C0",X"18",X"DE",X"3A",X"83",X"4C",X"D7",
		X"07",X"E6",X"1C",X"CD",X"07",X"23",X"71",X"EB",X"70",X"3E",X"04",X"84",X"67",X"36",X"19",X"EB",
		X"3E",X"04",X"84",X"67",X"36",X"03",X"C9",X"21",X"24",X"23",X"CD",X"52",X"21",X"56",X"23",X"5E",
		X"23",X"4E",X"23",X"46",X"6A",X"16",X"40",X"62",X"7B",X"FE",X"A0",X"30",X"01",X"14",X"7D",X"FE",
		X"A0",X"D0",X"24",X"C9",X"AC",X"CA",X"F2",X"B5",X"AB",X"EA",X"F9",X"B4",X"CA",X"0A",X"F7",X"B6",
		X"EA",X"0B",X"F7",X"B7",X"0A",X"EC",X"F3",X"B0",X"0B",X"CC",X"FA",X"B1",X"EC",X"AC",X"F8",X"B2",
		X"CC",X"AB",X"F8",X"B3",X"21",X"00",X"40",X"06",X"10",X"CD",X"66",X"23",X"2E",X"20",X"06",X"10",
		X"CD",X"66",X"23",X"21",X"5F",X"40",X"11",X"20",X"00",X"36",X"40",X"19",X"06",X"0B",X"3A",X"9B",
		X"41",X"77",X"19",X"10",X"FC",X"C9",X"36",X"40",X"23",X"10",X"FB",X"C9",X"21",X"16",X"4E",X"7E",
		X"B7",X"C0",X"3A",X"01",X"4E",X"FE",X"10",X"D8",X"36",X"FF",X"21",X"1C",X"4C",X"3A",X"20",X"4C",
		X"CB",X"57",X"28",X"01",X"23",X"34",X"CD",X"AC",X"21",X"3A",X"90",X"50",X"E6",X"C0",X"C9",X"3A",
		X"D0",X"50",X"E6",X"30",X"FE",X"30",X"C0",X"00",X"00",X"FF",X"32",X"03",X"4E",X"3A",X"06",X"4E",
		X"21",X"00",X"09",X"FE",X"08",X"30",X"11",X"B7",X"21",X"05",X"00",X"28",X"0B",X"47",X"7D",X"85",
		X"27",X"6F",X"7C",X"8C",X"27",X"67",X"10",X"F6",X"22",X"0E",X"4E",X"C9",X"3A",X"83",X"4C",X"47",
		X"E6",X"0F",X"C0",X"21",X"20",X"4C",X"7E",X"E6",X"07",X"28",X"16",X"CB",X"56",X"28",X"09",X"CB",
		X"60",X"20",X"0E",X"21",X"C5",X"43",X"18",X"1F",X"CB",X"60",X"20",X"05",X"21",X"D8",X"43",X"18",
		X"16",X"21",X"C5",X"43",X"36",X"50",X"23",X"36",X"55",X"23",X"36",X"02",X"2E",X"D8",X"36",X"50",
		X"23",X"36",X"55",X"23",X"36",X"01",X"C9",X"06",X"03",X"C3",X"66",X"23",X"3A",X"90",X"4C",X"B7",
		X"C8",X"21",X"10",X"40",X"06",X"10",X"FE",X"01",X"CA",X"66",X"23",X"3A",X"20",X"4C",X"CB",X"57",
		X"3A",X"1C",X"4C",X"28",X"03",X"3A",X"1D",X"4C",X"FE",X"02",X"D0",X"21",X"1D",X"40",X"11",X"35",
		X"24",X"06",X"0A",X"1A",X"77",X"2B",X"13",X"10",X"FA",X"06",X"0A",X"7C",X"C6",X"04",X"67",X"23",
		X"36",X"03",X"10",X"FB",X"C9",X"47",X"41",X"4D",X"45",X"40",X"4F",X"56",X"45",X"52",X"40",X"21",
		X"E4",X"4F",X"7E",X"23",X"B6",X"E6",X"07",X"2B",X"20",X"1D",X"E5",X"7D",X"D6",X"10",X"6F",X"7E",
		X"D7",X"E5",X"CD",X"CB",X"13",X"E1",X"E6",X"0F",X"47",X"A6",X"E6",X"0F",X"20",X"01",X"77",X"23",
		X"7E",X"2B",X"A0",X"28",X"01",X"77",X"E1",X"CD",X"48",X"2D",X"18",X"D6",X"21",X"80",X"4E",X"11",
		X"00",X"4F",X"01",X"80",X"00",X"ED",X"B0",X"CD",X"81",X"24",X"CD",X"4F",X"25",X"CD",X"0B",X"25",
		X"C9",X"21",X"60",X"40",X"11",X"80",X"4E",X"CD",X"74",X"21",X"30",X"12",X"47",X"CD",X"FD",X"24",
		X"78",X"20",X"0B",X"36",X"FF",X"CD",X"B5",X"24",X"7D",X"E6",X"1F",X"B0",X"12",X"13",X"23",X"7D",
		X"E6",X"1F",X"20",X"02",X"12",X"13",X"7D",X"FE",X"BF",X"20",X"DC",X"7C",X"FE",X"43",X"20",X"D7",
		X"AF",X"12",X"13",X"12",X"C9",X"E5",X"21",X"CD",X"24",X"06",X"00",X"BE",X"28",X"04",X"04",X"23",
		X"18",X"F9",X"78",X"07",X"07",X"07",X"07",X"07",X"E6",X"E0",X"47",X"E1",X"C9",X"A7",X"A7",X"A7",
		X"A7",X"A7",X"A7",X"A7",X"A7",X"A8",X"A9",X"A8",X"A9",X"A8",X"A9",X"A8",X"A9",X"AA",X"AB",X"AA",
		X"AB",X"AA",X"AB",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"BA",X"BB",X"BC",X"BD",X"B8",X"B9",X"B8",
		X"B9",X"B8",X"B9",X"B8",X"B9",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"E5",X"3E",X"04",
		X"84",X"67",X"7E",X"E1",X"CD",X"47",X"1D",X"C8",X"FE",X"03",X"C9",X"21",X"60",X"40",X"11",X"00",
		X"4F",X"4D",X"1A",X"B7",X"20",X"07",X"69",X"CD",X"50",X"21",X"4D",X"18",X"0D",X"E6",X"1F",X"47",
		X"7D",X"E6",X"E0",X"B0",X"6F",X"1A",X"CD",X"36",X"25",X"77",X"13",X"7C",X"FE",X"43",X"20",X"E2",
		X"7D",X"FE",X"BF",X"38",X"DD",X"C9",X"E5",X"0F",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",X"47",X"CD",
		X"00",X"20",X"87",X"87",X"87",X"B0",X"21",X"CD",X"24",X"CD",X"52",X"21",X"7E",X"E1",X"C9",X"21",
		X"40",X"40",X"11",X"40",X"44",X"1A",X"F5",X"7E",X"E5",X"21",X"8D",X"25",X"CD",X"84",X"25",X"E1",
		X"20",X"09",X"CD",X"9B",X"25",X"1A",X"E6",X"1F",X"B0",X"18",X"03",X"1A",X"E6",X"1F",X"12",X"F1",
		X"E6",X"E0",X"28",X"03",X"CD",X"C9",X"25",X"23",X"13",X"7D",X"FE",X"BF",X"20",X"D7",X"7C",X"FE",
		X"43",X"20",X"D2",X"C9",X"46",X"23",X"BE",X"23",X"C8",X"10",X"FB",X"04",X"C9",X"0D",X"FF",X"D2",
		X"FC",X"FE",X"FD",X"D1",X"E1",X"E5",X"EA",X"CC",X"CD",X"CE",X"CF",X"06",X"E0",X"D6",X"CC",X"28",
		X"25",X"06",X"C0",X"3D",X"28",X"20",X"06",X"A0",X"3D",X"28",X"1B",X"06",X"80",X"3D",X"28",X"16",
		X"1A",X"E6",X"1F",X"06",X"60",X"FE",X"06",X"C8",X"FE",X"02",X"C8",X"FE",X"04",X"C8",X"06",X"40",
		X"FE",X"03",X"C8",X"06",X"00",X"C9",X"36",X"FF",X"C9",X"D7",X"0F",X"E6",X"07",X"47",X"05",X"05",
		X"28",X"18",X"05",X"28",X"0F",X"0E",X"CF",X"05",X"28",X"09",X"0D",X"05",X"28",X"05",X"0D",X"05",
		X"28",X"01",X"0D",X"71",X"1A",X"CD",X"6D",X"1D",X"12",X"C9",X"1A",X"E6",X"E0",X"F6",X"03",X"12",
		X"C9",X"21",X"14",X"4E",X"3A",X"E7",X"41",X"FE",X"D8",X"28",X"0A",X"CB",X"8E",X"21",X"F0",X"41",
		X"CD",X"2E",X"2F",X"18",X"08",X"CB",X"CE",X"21",X"E7",X"41",X"CD",X"2E",X"2F",X"21",X"14",X"4E",
		X"3A",X"74",X"41",X"FE",X"DC",X"28",X"08",X"CB",X"86",X"21",X"94",X"42",X"C3",X"28",X"2F",X"CB",
		X"C6",X"21",X"74",X"41",X"C3",X"28",X"2F",X"3A",X"14",X"4E",X"0F",X"38",X"05",X"CD",X"DA",X"2E",
		X"18",X"03",X"CD",X"E2",X"2E",X"3A",X"14",X"4E",X"0F",X"0F",X"DA",X"FA",X"2E",X"C3",X"F2",X"2E",
		X"3A",X"11",X"4E",X"B7",X"20",X"0C",X"11",X"CE",X"4F",X"21",X"E4",X"4F",X"01",X"A8",X"4C",X"CD",
		X"79",X"26",X"11",X"92",X"4C",X"21",X"E8",X"4F",X"01",X"A9",X"4C",X"CD",X"79",X"26",X"11",X"94",
		X"4C",X"21",X"EA",X"4F",X"01",X"AA",X"4C",X"CD",X"79",X"26",X"3A",X"07",X"4E",X"E6",X"81",X"E8",
		X"11",X"96",X"4C",X"21",X"EC",X"4F",X"01",X"AB",X"4C",X"1A",X"07",X"30",X"0C",X"E5",X"CD",X"3F",
		X"2C",X"E1",X"7E",X"23",X"B6",X"E6",X"07",X"C8",X"2B",X"E5",X"CD",X"92",X"26",X"E1",X"C8",X"C3",
		X"3F",X"2C",X"1A",X"E6",X"0F",X"87",X"21",X"B4",X"26",X"CD",X"52",X"21",X"0A",X"3C",X"FE",X"10",
		X"38",X"01",X"AF",X"02",X"47",X"04",X"AF",X"4F",X"37",X"17",X"CB",X"11",X"10",X"FB",X"A6",X"C0",
		X"79",X"23",X"A6",X"C9",X"00",X"80",X"80",X"80",X"20",X"84",X"88",X"88",X"48",X"92",X"92",X"92",
		X"2A",X"95",X"AA",X"AA",X"5A",X"DA",X"6D",X"6D",X"6D",X"DB",X"77",X"77",X"DE",X"F7",X"7F",X"7F",
		X"7F",X"FF",X"FF",X"FF",X"00",X"59",X"AA",X"00",X"00",X"EF",X"25",X"04",X"0C",X"0B",X"00",X"B2",
		X"7D",X"00",X"00",X"97",X"23",X"04",X"05",X"07",X"00",X"B0",X"CE",X"00",X"00",X"81",X"25",X"04",
		X"05",X"17",X"00",X"B3",X"6D",X"00",X"00",X"E9",X"26",X"04",X"05",X"0F",X"00",X"B0",X"D4",X"00",
		X"00",X"49",X"26",X"04",X"05",X"1F",X"00",X"B2",X"7D",X"AF",X"00",X"DF",X"26",X"14",X"0E",X"CB",
		X"00",X"B0",X"CE",X"AF",X"00",X"F3",X"26",X"14",X"0E",X"CB",X"10",X"B3",X"6D",X"AF",X"00",X"11",
		X"27",X"14",X"0E",X"CB",X"08",X"B0",X"D4",X"AF",X"00",X"FD",X"26",X"14",X"0E",X"CB",X"18",X"B8",
		X"BB",X"AF",X"00",X"7B",X"26",X"14",X"0E",X"CB",X"20",X"B9",X"AB",X"AF",X"00",X"CD",X"24",X"14",
		X"0E",X"CB",X"28",X"B9",X"B6",X"AF",X"00",X"07",X"27",X"14",X"0E",X"CB",X"38",X"B2",X"7E",X"00",
		X"00",X"E1",X"24",X"14",X"06",X"ED",X"6F",X"B3",X"6E",X"00",X"00",X"17",X"26",X"14",X"06",X"ED",
		X"67",X"4E",X"16",X"00",X"00",X"CB",X"26",X"14",X"0F",X"CB",X"40",X"B7",X"B6",X"00",X"00",X"8F",
		X"26",X"14",X"0F",X"CB",X"C0",X"B1",X"75",X"00",X"00",X"25",X"27",X"14",X"0F",X"CB",X"80",X"80",
		X"B2",X"00",X"00",X"39",X"27",X"04",X"09",X"C3",X"00",X"80",X"E4",X"00",X"00",X"75",X"27",X"04",
		X"09",X"C2",X"00",X"82",X"A0",X"00",X"00",X"67",X"26",X"04",X"09",X"CA",X"00",X"80",X"CD",X"00",
		X"00",X"2D",X"24",X"04",X"09",X"D2",X"00",X"7F",X"08",X"00",X"00",X"2B",X"26",X"04",X"09",X"DA",
		X"00",X"81",X"29",X"00",X"00",X"AD",X"26",X"04",X"09",X"E2",X"00",X"81",X"1F",X"00",X"00",X"1B",
		X"27",X"04",X"09",X"EA",X"00",X"81",X"10",X"00",X"00",X"3F",X"26",X"04",X"09",X"F2",X"00",X"80",
		X"98",X"00",X"00",X"61",X"27",X"04",X"09",X"FA",X"00",X"80",X"D9",X"00",X"00",X"00",X"00",X"14",
		X"09",X"E2",X"00",X"80",X"E8",X"00",X"00",X"B1",X"27",X"14",X"09",X"EA",X"00",X"80",X"B2",X"AF",
		X"00",X"7F",X"27",X"14",X"10",X"18",X"00",X"81",X"6D",X"00",X"00",X"4D",X"27",X"14",X"10",X"D9",
		X"21",X"83",X"4C",X"7E",X"E6",X"FE",X"FE",X"4E",X"20",X"0B",X"7E",X"2F",X"32",X"07",X"50",X"0F",
		X"38",X"03",X"CD",X"00",X"18",X"21",X"1E",X"4C",X"11",X"36",X"40",X"01",X"00",X"01",X"CD",X"61",
		X"28",X"21",X"80",X"4C",X"11",X"F3",X"43",X"CD",X"58",X"28",X"3A",X"87",X"4C",X"B7",X"21",X"00",
		X"4E",X"3A",X"20",X"4C",X"E6",X"03",X"20",X"03",X"21",X"00",X"4D",X"3A",X"20",X"4C",X"CB",X"57",
		X"20",X"0C",X"1E",X"FD",X"CD",X"58",X"28",X"21",X"80",X"4D",X"1E",X"E8",X"18",X"0A",X"1E",X"E8",
		X"CD",X"58",X"28",X"21",X"00",X"4D",X"1E",X"FD",X"01",X"FF",X"03",X"CD",X"61",X"28",X"AF",X"12",
		X"C9",X"7E",X"D7",X"CD",X"6E",X"28",X"7E",X"CD",X"6E",X"28",X"23",X"10",X"F4",X"C9",X"E6",X"0F",
		X"CB",X"09",X"30",X"09",X"B7",X"28",X"04",X"0E",X"00",X"18",X"02",X"3E",X"40",X"12",X"1B",X"C9",
		X"E1",X"46",X"23",X"5E",X"23",X"56",X"23",X"EB",X"1A",X"77",X"D5",X"11",X"20",X"00",X"19",X"D1",
		X"13",X"10",X"F5",X"EB",X"E9",X"08",X"7B",X"D6",X"20",X"ED",X"44",X"47",X"08",X"77",X"3C",X"23",
		X"10",X"FB",X"19",X"0D",X"20",X"EF",X"C9",X"08",X"7B",X"D6",X"20",X"ED",X"44",X"47",X"08",X"77",
		X"23",X"10",X"FC",X"19",X"0D",X"20",X"F0",X"C9",X"21",X"76",X"42",X"11",X"1D",X"00",X"3E",X"0A",
		X"0E",X"03",X"CD",X"95",X"28",X"21",X"76",X"46",X"3E",X"1D",X"0E",X"03",X"CD",X"A7",X"28",X"3E",
		X"1F",X"32",X"78",X"46",X"32",X"98",X"46",X"32",X"B8",X"46",X"C9",X"3E",X"13",X"32",X"97",X"42",
		X"3C",X"32",X"B7",X"42",X"C9",X"21",X"76",X"42",X"11",X"1E",X"00",X"3E",X"40",X"0E",X"03",X"CD",
		X"A7",X"28",X"3E",X"EE",X"32",X"76",X"42",X"32",X"96",X"42",X"3E",X"F7",X"32",X"B6",X"42",X"3E",
		X"1E",X"32",X"B8",X"46",X"3E",X"03",X"32",X"76",X"46",X"32",X"96",X"46",X"32",X"B6",X"46",X"C9",
		X"21",X"D6",X"40",X"11",X"1D",X"00",X"3E",X"16",X"0E",X"03",X"CD",X"95",X"28",X"21",X"D6",X"44",
		X"3E",X"09",X"0E",X"03",X"C3",X"A7",X"28",X"21",X"D7",X"40",X"11",X"1E",X"00",X"3E",X"1F",X"0E",
		X"03",X"C3",X"95",X"28",X"21",X"D7",X"40",X"11",X"1E",X"00",X"3E",X"40",X"0E",X"03",X"CD",X"A7",
		X"28",X"21",X"D8",X"40",X"36",X"F8",X"2E",X"F8",X"36",X"F8",X"21",X"17",X"41",X"36",X"FA",X"23",
		X"36",X"F4",X"3E",X"03",X"21",X"D8",X"44",X"77",X"2E",X"F8",X"77",X"21",X"17",X"45",X"77",X"23",
		X"77",X"C9",X"21",X"E3",X"42",X"11",X"1C",X"00",X"3E",X"25",X"0E",X"04",X"CD",X"95",X"28",X"2E",
		X"43",X"36",X"F3",X"2E",X"47",X"77",X"2E",X"27",X"36",X"31",X"3E",X"1C",X"21",X"E3",X"46",X"1B",
		X"0E",X"04",X"CD",X"A7",X"28",X"3E",X"03",X"21",X"E7",X"46",X"77",X"21",X"07",X"47",X"77",X"2E",
		X"43",X"77",X"2E",X"04",X"36",X"0F",X"23",X"36",X"14",X"3E",X"1D",X"32",X"E5",X"46",X"C9",X"21",
		X"04",X"43",X"36",X"36",X"23",X"36",X"37",X"C9",X"3E",X"F9",X"32",X"E5",X"42",X"21",X"04",X"43",
		X"36",X"36",X"23",X"36",X"40",X"C9",X"21",X"50",X"40",X"36",X"5C",X"23",X"36",X"5D",X"23",X"36",
		X"5E",X"21",X"6F",X"40",X"11",X"1C",X"00",X"3E",X"5F",X"0E",X"03",X"CD",X"95",X"28",X"23",X"77",
		X"23",X"3C",X"77",X"23",X"3C",X"77",X"21",X"4F",X"44",X"3E",X"0D",X"0E",X"05",X"CD",X"A7",X"28",
		X"21",X"6F",X"44",X"3E",X"0B",X"77",X"2E",X"8F",X"77",X"23",X"36",X"0C",X"C9",X"21",X"51",X"40",
		X"11",X"1E",X"00",X"3E",X"6E",X"0E",X"02",X"CD",X"95",X"28",X"21",X"B1",X"40",X"3E",X"72",X"0E",
		X"02",X"C3",X"95",X"28",X"21",X"6F",X"40",X"11",X"1E",X"00",X"3E",X"7E",X"0E",X"02",X"CD",X"95",
		X"28",X"21",X"51",X"40",X"36",X"5D",X"23",X"36",X"5E",X"19",X"23",X"36",X"61",X"23",X"36",X"62",
		X"21",X"B1",X"40",X"3E",X"76",X"0E",X"02",X"C3",X"95",X"28",X"3E",X"82",X"32",X"8F",X"40",X"21",
		X"51",X"40",X"3E",X"6E",X"11",X"1E",X"00",X"0E",X"02",X"CD",X"95",X"28",X"21",X"B1",X"40",X"3E",
		X"7A",X"0E",X"02",X"C3",X"95",X"28",X"21",X"3B",X"43",X"11",X"1C",X"00",X"0E",X"03",X"3E",X"83",
		X"CD",X"95",X"28",X"21",X"3B",X"47",X"0E",X"03",X"3E",X"1B",X"C3",X"A7",X"28",X"21",X"3C",X"43",
		X"36",X"8F",X"23",X"36",X"90",X"C9",X"21",X"3B",X"43",X"11",X"1C",X"00",X"0E",X"03",X"3E",X"95",
		X"CD",X"95",X"28",X"21",X"3B",X"47",X"0E",X"03",X"3E",X"09",X"C3",X"A7",X"28",X"21",X"3D",X"43",
		X"11",X"1E",X"00",X"3E",X"A1",X"0E",X"03",X"CD",X"95",X"28",X"21",X"5C",X"43",X"36",X"A3",X"23",
		X"36",X"9B",X"C9",X"11",X"80",X"4C",X"21",X"00",X"4E",X"06",X"03",X"1A",X"BE",X"20",X"05",X"23",
		X"13",X"10",X"F8",X"C9",X"D0",X"2E",X"00",X"1E",X"80",X"01",X"03",X"00",X"ED",X"B0",X"3A",X"40",
		X"50",X"0F",X"0F",X"C9",X"3A",X"83",X"4C",X"FE",X"A9",X"C0",X"CD",X"D0",X"3A",X"C8",X"00",X"00",
		X"ED",X"B0",X"C9",X"7E",X"81",X"77",X"FE",X"04",X"D8",X"D6",X"04",X"77",X"06",X"02",X"CD",X"DA",
		X"2A",X"06",X"03",X"CD",X"DA",X"2A",X"CD",X"C0",X"31",X"C9",X"37",X"2B",X"7E",X"CE",X"00",X"27",
		X"77",X"10",X"F8",X"C9",X"21",X"D4",X"4F",X"46",X"21",X"C4",X"4F",X"4E",X"78",X"E6",X"0F",X"C8",
		X"78",X"0F",X"30",X"06",X"CB",X"D9",X"CB",X"81",X"18",X"19",X"0F",X"30",X"06",X"CB",X"99",X"CB",
		X"C9",X"18",X"10",X"0F",X"30",X"06",X"CB",X"99",X"CB",X"89",X"18",X"07",X"0F",X"30",X"04",X"CB",
		X"D9",X"CB",X"C1",X"71",X"11",X"8F",X"4C",X"1A",X"3C",X"12",X"4F",X"78",X"E6",X"09",X"20",X"3D",
		X"78",X"E6",X"06",X"20",X"08",X"3A",X"D5",X"4F",X"47",X"E6",X"09",X"20",X"30",X"79",X"FE",X"04",
		X"20",X"05",X"CB",X"D6",X"CB",X"86",X"C9",X"FE",X"08",X"20",X"05",X"CB",X"D6",X"CB",X"C6",X"C9",
		X"FE",X"0C",X"20",X"04",X"CB",X"96",X"18",X"F5",X"FE",X"10",X"20",X"02",X"18",X"ED",X"FE",X"14",
		X"20",X"02",X"18",X"DE",X"FE",X"18",X"C0",X"CB",X"96",X"CB",X"86",X"18",X"2F",X"79",X"FE",X"04",
		X"20",X"05",X"CB",X"D6",X"CB",X"8E",X"C9",X"FE",X"08",X"20",X"05",X"CB",X"D6",X"CB",X"CE",X"C9",
		X"FE",X"0C",X"20",X"05",X"CB",X"96",X"CB",X"CE",X"C9",X"FE",X"10",X"20",X"02",X"18",X"EC",X"FE",
		X"14",X"20",X"02",X"18",X"DD",X"FE",X"18",X"C0",X"CB",X"96",X"CB",X"8E",X"AF",X"12",X"C9",X"E5",
		X"D5",X"CD",X"51",X"3A",X"D1",X"E1",X"3E",X"7F",X"20",X"02",X"1A",X"96",X"13",X"23",X"F0",X"ED",
		X"44",X"C9",X"CD",X"8F",X"2B",X"4F",X"18",X"F2",X"3A",X"11",X"4E",X"B7",X"C0",X"21",X"E8",X"4F",
		X"06",X"02",X"11",X"E4",X"4F",X"CD",X"A2",X"2B",X"81",X"38",X"05",X"FE",X"08",X"DC",X"C3",X"2B",
		X"10",X"F0",X"C9",X"E5",X"7D",X"D6",X"22",X"6F",X"CB",X"5E",X"E1",X"C0",X"3E",X"83",X"32",X"5C",
		X"4C",X"3E",X"FF",X"32",X"90",X"4C",X"21",X"20",X"4C",X"CB",X"F6",X"F1",X"C9",X"11",X"1E",X"4C",
		X"CD",X"23",X"2C",X"21",X"20",X"4C",X"7E",X"0F",X"D8",X"0F",X"D8",X"1A",X"B7",X"C8",X"FE",X"01",
		X"3A",X"01",X"4C",X"4F",X"3A",X"40",X"50",X"28",X"1C",X"CB",X"77",X"20",X"18",X"36",X"83",X"1A",
		X"3D",X"3D",X"27",X"12",X"21",X"1C",X"4C",X"71",X"23",X"71",X"AF",X"32",X"87",X"4C",X"32",X"90",
		X"4C",X"32",X"5C",X"4C",X"C9",X"CB",X"6F",X"C0",X"36",X"81",X"1A",X"3D",X"27",X"12",X"21",X"1C",
		X"4C",X"18",X"E6",X"21",X"83",X"4C",X"7E",X"E6",X"FE",X"FE",X"08",X"C0",X"7E",X"2F",X"32",X"07",
		X"50",X"0F",X"D8",X"C3",X"B5",X"3A",X"EB",X"35",X"EB",X"C0",X"13",X"1A",X"1B",X"12",X"C9",X"E5",
		X"7D",X"D6",X"10",X"6F",X"7E",X"0F",X"E1",X"23",X"30",X"01",X"34",X"2B",X"0F",X"30",X"01",X"34",
		X"0F",X"30",X"01",X"35",X"0F",X"D0",X"23",X"35",X"2B",X"C9",X"CD",X"E9",X"2D",X"0C",X"C2",X"4F",
		X"B4",X"83",X"F8",X"01",X"00",X"83",X"48",X"09",X"48",X"09",X"00",X"00",X"CD",X"E9",X"2D",X"0C",
		X"E2",X"4F",X"00",X"00",X"88",X"18",X"00",X"00",X"A0",X"B0",X"70",X"B0",X"01",X"01",X"C9",X"7E",
		X"D6",X"10",X"0F",X"0F",X"0F",X"E6",X"1F",X"57",X"23",X"7E",X"2B",X"D6",X"10",X"2F",X"06",X"03",
		X"CB",X"3A",X"1F",X"10",X"FB",X"5F",X"C9",X"21",X"8C",X"4C",X"7E",X"3C",X"77",X"FE",X"08",X"D8",
		X"36",X"00",X"21",X"D8",X"4F",X"CD",X"C0",X"2C",X"23",X"23",X"7D",X"FE",X"DC",X"20",X"F6",X"3A",
		X"10",X"4E",X"B7",X"C8",X"CD",X"00",X"20",X"3D",X"28",X"2B",X"3D",X"28",X"19",X"3D",X"28",X"16",
		X"E5",X"46",X"7D",X"D6",X"10",X"6F",X"4E",X"78",X"E6",X"06",X"79",X"20",X"04",X"EE",X"02",X"18",
		X"02",X"EE",X"01",X"77",X"E1",X"C9",X"3A",X"07",X"4E",X"E6",X"81",X"E8",X"7D",X"D6",X"10",X"6F",
		X"7E",X"EE",X"04",X"77",X"C9",X"21",X"CC",X"4F",X"7E",X"E6",X"FC",X"77",X"C9",X"21",X"D8",X"4F",
		X"46",X"7D",X"D6",X"10",X"6F",X"7E",X"CB",X"08",X"30",X"06",X"CB",X"D7",X"CB",X"87",X"18",X"18",
		X"CB",X"08",X"30",X"06",X"CB",X"97",X"CB",X"CF",X"18",X"0E",X"CB",X"08",X"30",X"04",X"E6",X"F9",
		X"18",X"06",X"CB",X"08",X"30",X"02",X"F6",X"05",X"77",X"7D",X"C6",X"12",X"6F",X"FE",X"DC",X"28",
		X"05",X"FE",X"DE",X"38",X"CB",X"C9",X"3A",X"10",X"4E",X"B7",X"C8",X"CD",X"00",X"20",X"FE",X"02",
		X"28",X"05",X"FE",X"03",X"C8",X"18",X"B9",X"46",X"21",X"CC",X"4F",X"CB",X"48",X"20",X"06",X"CB",
		X"50",X"C8",X"CB",X"8E",X"C9",X"CB",X"CE",X"C9",X"23",X"23",X"7D",X"FE",X"E6",X"28",X"F9",X"FE",
		X"EE",X"D8",X"33",X"33",X"C9",X"21",X"E8",X"4F",X"06",X"02",X"11",X"E6",X"4F",X"CD",X"61",X"3A",
		X"81",X"38",X"05",X"FE",X"05",X"DC",X"6B",X"2D",X"10",X"F0",X"C9",X"3A",X"C6",X"4F",X"E6",X"F8",
		X"FE",X"B8",X"C0",X"E5",X"7D",X"FE",X"EA",X"3E",X"FF",X"21",X"CA",X"4F",X"28",X"09",X"CB",X"5E",
		X"20",X"1D",X"32",X"EF",X"4F",X"18",X"09",X"2B",X"2B",X"CB",X"5E",X"20",X"12",X"32",X"EE",X"4F",
		X"CB",X"DE",X"23",X"36",X"10",X"CD",X"EE",X"31",X"CD",X"57",X"2F",X"21",X"1B",X"4E",X"34",X"E1",
		X"C9",X"21",X"00",X"4D",X"11",X"00",X"4E",X"18",X"16",X"21",X"80",X"4D",X"11",X"00",X"4E",X"18",
		X"0E",X"21",X"00",X"4E",X"11",X"00",X"4D",X"18",X"06",X"21",X"00",X"4E",X"11",X"80",X"4D",X"01",
		X"40",X"00",X"ED",X"B0",X"C9",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"77",X"23",X"0D",X"20",X"FB",
		X"C9",X"CD",X"CB",X"2D",X"10",X"FB",X"C9",X"AF",X"18",X"02",X"3E",X"01",X"32",X"03",X"50",X"C9",
		X"AF",X"18",X"02",X"3E",X"01",X"32",X"01",X"50",X"C9",X"E1",X"46",X"23",X"5E",X"23",X"56",X"23",
		X"7E",X"23",X"12",X"13",X"10",X"FA",X"E9",X"3A",X"20",X"4C",X"47",X"E6",X"03",X"28",X"18",X"CB",
		X"50",X"3A",X"00",X"50",X"28",X"07",X"CB",X"67",X"28",X"03",X"3A",X"40",X"50",X"32",X"8D",X"4C",
		X"CD",X"37",X"2F",X"79",X"32",X"D5",X"4F",X"21",X"83",X"4C",X"7E",X"E6",X"0E",X"FE",X"02",X"C0",
		X"7E",X"2F",X"32",X"07",X"50",X"0F",X"D8",X"C3",X"00",X"18",X"CD",X"E9",X"2D",X"06",X"38",X"40",
		X"54",X"49",X"44",X"45",X"52",X"43",X"CD",X"4C",X"2E",X"CD",X"E9",X"2D",X"03",X"D8",X"43",X"50",
		X"55",X"01",X"CD",X"E9",X"2D",X"03",X"C5",X"43",X"50",X"55",X"02",X"C9",X"CD",X"E9",X"2D",X"08",
		X"CC",X"43",X"45",X"52",X"4F",X"43",X"53",X"40",X"49",X"48",X"C9",X"21",X"00",X"44",X"01",X"00",
		X"04",X"CD",X"D1",X"2D",X"C9",X"21",X"00",X"40",X"01",X"00",X"04",X"CD",X"D1",X"2D",X"C9",X"21",
		X"00",X"30",X"11",X"40",X"40",X"01",X"C0",X"02",X"7E",X"D7",X"F6",X"F0",X"12",X"13",X"7E",X"F6",
		X"F0",X"12",X"13",X"23",X"0D",X"20",X"F1",X"10",X"EF",X"CD",X"E9",X"2D",X"0A",X"C7",X"41",X"E0",
		X"E1",X"E1",X"E2",X"D3",X"E3",X"E1",X"E1",X"E2",X"E3",X"CD",X"E9",X"2D",X"0A",X"27",X"42",X"E4",
		X"E5",X"E5",X"E6",X"E5",X"E7",X"E5",X"E5",X"E6",X"E7",X"3E",X"D2",X"32",X"48",X"40",X"32",X"54",
		X"40",X"32",X"61",X"40",X"32",X"E0",X"41",X"CD",X"F2",X"2E",X"CD",X"80",X"28",X"0A",X"73",X"41",
		X"E8",X"E8",X"E8",X"E9",X"EA",X"EA",X"EB",X"E8",X"E8",X"EC",X"CD",X"80",X"28",X"0A",X"76",X"41",
		X"ED",X"EE",X"EE",X"EF",X"D1",X"D1",X"ED",X"EE",X"EE",X"EE",X"21",X"94",X"42",X"11",X"DF",X"DE",
		X"18",X"06",X"21",X"74",X"41",X"11",X"DD",X"DC",X"CD",X"0F",X"2F",X"72",X"23",X"CD",X"0F",X"2F",
		X"73",X"C9",X"21",X"F0",X"41",X"11",X"DB",X"DA",X"18",X"06",X"21",X"E7",X"41",X"11",X"D9",X"D8",
		X"CD",X"0F",X"2F",X"72",X"D5",X"11",X"20",X"00",X"19",X"D1",X"CD",X"0F",X"2F",X"73",X"C9",X"7E",
		X"CD",X"1F",X"2F",X"C0",X"E5",X"21",X"05",X"4E",X"0E",X"01",X"CD",X"C3",X"2A",X"E1",X"C9",X"D6",
		X"CC",X"C8",X"3D",X"C8",X"3D",X"C8",X"3D",X"C9",X"36",X"FF",X"23",X"36",X"FF",X"C9",X"36",X"FF",
		X"11",X"20",X"00",X"19",X"36",X"FF",X"C9",X"06",X"04",X"0E",X"01",X"0F",X"D0",X"CB",X"21",X"10",
		X"FA",X"C9",X"21",X"40",X"44",X"7E",X"E6",X"E0",X"F6",X"03",X"77",X"23",X"7C",X"FE",X"47",X"20",
		X"F4",X"7D",X"FE",X"C0",X"C8",X"18",X"EE",X"2A",X"0E",X"4E",X"7C",X"FE",X"10",X"38",X"03",X"21",
		X"00",X"09",X"11",X"02",X"4E",X"CD",X"29",X"3A",X"E5",X"CD",X"39",X"3A",X"22",X"0E",X"4E",X"E1",
		X"CD",X"F7",X"39",X"2A",X"C4",X"4F",X"E5",X"2A",X"C6",X"4F",X"E5",X"AF",X"32",X"C7",X"4F",X"ED",
		X"53",X"C4",X"4F",X"3A",X"83",X"4C",X"C6",X"60",X"47",X"3A",X"83",X"4C",X"B8",X"20",X"FA",X"E1",
		X"22",X"C6",X"4F",X"E1",X"22",X"C4",X"4F",X"C9",X"00",X"8B",X"2F",X"15",X"00",X"FE",X"4E",X"B9",
		X"FB",X"83",X"D5",X"95",X"2F",X"15",X"00",X"00",X"4F",X"B9",X"FB",X"83",X"C7",X"9F",X"2F",X"15",
		X"00",X"7E",X"4F",X"B2",X"81",X"A7",X"30",X"6D",X"2F",X"15",X"00",X"14",X"4E",X"92",X"CE",X"7A",
		X"C0",X"79",X"28",X"15",X"00",X"16",X"4E",X"A6",X"13",X"56",X"36",X"27",X"2F",X"15",X"00",X"1C",
		X"4C",X"A6",X"13",X"14",X"E7",X"C7",X"2F",X"15",X"00",X"1D",X"4C",X"92",X"30",X"5C",X"A8",X"A9",
		X"2F",X"15",X"00",X"9F",X"4C",X"B0",X"CB",X"98",X"08",X"55",X"2E",X"15",X"00",X"A0",X"4C",X"59",
		X"EF",X"9E",X"D6",X"B9",X"2E",X"15",X"00",X"A2",X"4C",X"5C",X"4E",X"4E",X"91",X"31",X"2F",X"EF",
		X"0A",X"AA",X"AA",X"A4",X"FC",X"3A",X"AA",X"A0",X"00",X"08",X"FC",X"3A",X"AA",X"AA",X"AA",X"A0",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",X"00",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"C7",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"00",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"8F",X"F1",X"2F",X"F5",X"FF",X"19",X"2F",X"F7",X"00",X"08",X"FF",X"19",X"2F",X"F1",X"2F",X"F7",
		X"8F",X"F7",X"8F",X"FB",X"FF",X"70",X"8F",X"F3",X"AA",X"A4",X"FF",X"70",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"F7",X"8F",X"FB",X"FF",X"70",X"8F",X"FF",X"FF",X"FF",X"FF",X"70",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"F3",X"4F",X"F6",X"FF",X"3A",X"4F",X"FF",X"FF",X"FF",X"FF",X"3A",X"4F",X"F3",X"4F",X"F7",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F1",X"2F",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F3",X"4F",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"8F",X"F1",X"2F",X"F5",X"FF",X"19",X"2F",X"FF",X"FF",X"F0",X"FF",X"09",X"2F",X"F1",X"2F",X"F7",
		X"8F",X"F7",X"8F",X"FB",X"FF",X"70",X"8F",X"FF",X"FF",X"F0",X"FF",X"00",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"F7",X"8F",X"FB",X"FF",X"70",X"8F",X"F1",X"2F",X"F0",X"FF",X"00",X"8F",X"F7",X"8F",X"F7",
		X"4F",X"F3",X"4F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F0",X"FF",X"0A",X"4F",X"F3",X"4F",X"F3",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"0F",X"FF",X"FF",X"FF",X"FC",
		X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"0F",X"FF",X"FF",X"FF",X"FD",
		X"2F",X"F1",X"2F",X"F0",X"00",X"00",X"00",X"00",X"0F",X"F0",X"FF",X"09",X"2F",X"F1",X"2F",X"F1",
		X"8F",X"F7",X"8F",X"FB",X"FF",X"70",X"8F",X"F7",X"8F",X"F0",X"FF",X"00",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"F7",X"8F",X"FB",X"FF",X"70",X"8F",X"F7",X"8F",X"F0",X"FF",X"00",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"F3",X"4F",X"F6",X"FF",X"3A",X"4F",X"F3",X"4F",X"F0",X"FF",X"00",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"70",X"8F",X"F7",X"8F",X"F7",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"4F",X"F3",X"4F",X"F7",
		X"8F",X"F1",X"99",X"92",X"FF",X"19",X"2F",X"F1",X"2F",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",
		X"8F",X"F7",X"00",X"08",X"FF",X"3A",X"4F",X"F7",X"8F",X"FB",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",
		X"8F",X"F7",X"00",X"08",X"FF",X"FF",X"FF",X"F7",X"8F",X"FB",X"FF",X"19",X"2F",X"F1",X"99",X"90",
		X"8F",X"F3",X"AA",X"A4",X"FF",X"FF",X"FF",X"F3",X"4F",X"F6",X"FF",X"3A",X"4F",X"F7",X"00",X"00",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"19",X"2F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"00",X"00",
		X"8E",X"FF",X"FF",X"FF",X"FF",X"70",X"8E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"D7",X"00",X"00",
		X"09",X"99",X"99",X"92",X"ED",X"70",X"09",X"99",X"99",X"92",X"ED",X"19",X"99",X"90",X"00",X"00",
		X"21",X"5E",X"4C",X"CB",X"46",X"C0",X"36",X"82",X"C9",X"21",X"5E",X"4C",X"36",X"81",X"C9",X"00",
		X"00",X"21",X"5E",X"4C",X"36",X"00",X"C9",X"21",X"5D",X"4C",X"7E",X"B7",X"C0",X"36",X"82",X"C9",
		X"21",X"5D",X"4C",X"36",X"00",X"23",X"23",X"36",X"81",X"C9",X"00",X"00",X"00",X"00",X"21",X"5D",
		X"4C",X"36",X"81",X"C9",X"21",X"5D",X"4C",X"36",X"85",X"C9",X"21",X"83",X"4C",X"7E",X"E6",X"FE",
		X"FE",X"A8",X"C0",X"7E",X"2F",X"32",X"07",X"50",X"0F",X"D8",X"C3",X"00",X"18",X"CD",X"FA",X"31",
		X"3A",X"20",X"4C",X"E6",X"03",X"C8",X"21",X"5C",X"4C",X"7E",X"B7",X"28",X"05",X"CD",X"82",X"32",
		X"18",X"5D",X"21",X"5D",X"4C",X"7E",X"23",X"23",X"B6",X"06",X"05",X"21",X"41",X"4C",X"CC",X"C5",
		X"2D",X"21",X"5D",X"4C",X"7E",X"23",X"B6",X"21",X"46",X"4C",X"06",X"05",X"CC",X"C5",X"2D",X"21",
		X"5E",X"4C",X"7E",X"B7",X"21",X"4B",X"4C",X"06",X"05",X"CC",X"C5",X"2D",X"21",X"5F",X"4C",X"7E",
		X"B7",X"C4",X"14",X"34",X"21",X"5E",X"4C",X"7E",X"CB",X"47",X"20",X"04",X"B7",X"C4",X"E1",X"33",
		X"21",X"5D",X"4C",X"7E",X"CB",X"47",X"20",X"05",X"CB",X"4F",X"C4",X"EC",X"33",X"21",X"5E",X"4C",
		X"7E",X"CB",X"47",X"C4",X"F7",X"33",X"21",X"5D",X"4C",X"7E",X"CB",X"47",X"C4",X"02",X"34",X"C3",
		X"08",X"33",X"CB",X"7F",X"CA",X"87",X"33",X"CB",X"BE",X"7E",X"E6",X"03",X"3D",X"21",X"9D",X"32",
		X"28",X"2F",X"3D",X"21",X"A9",X"32",X"28",X"29",X"21",X"B5",X"32",X"18",X"24",X"01",X"01",X"00",
		X"04",X"21",X"03",X"02",X"01",X"00",X"00",X"18",X"35",X"00",X"02",X"00",X"00",X"25",X"00",X"03",
		X"04",X"00",X"00",X"96",X"35",X"00",X"02",X"00",X"00",X"25",X"00",X"02",X"04",X"00",X"00",X"CA",
		X"35",X"11",X"50",X"4C",X"01",X"0C",X"00",X"ED",X"B0",X"CD",X"E3",X"2D",X"21",X"40",X"4C",X"06",
		X"10",X"C3",X"C5",X"2D",X"AF",X"32",X"58",X"4C",X"2A",X"5A",X"4C",X"7E",X"B7",X"CA",X"14",X"33",
		X"CD",X"19",X"33",X"3A",X"54",X"4C",X"CD",X"31",X"33",X"3A",X"50",X"4C",X"B7",X"28",X"14",X"23",
		X"3A",X"53",X"4C",X"CD",X"31",X"33",X"3A",X"50",X"4C",X"3D",X"28",X"07",X"23",X"3A",X"52",X"4C",
		X"CD",X"31",X"33",X"23",X"22",X"5A",X"4C",X"C9",X"21",X"40",X"4C",X"11",X"50",X"50",X"01",X"10",
		X"00",X"ED",X"B0",X"C9",X"11",X"D4",X"32",X"D5",X"E9",X"7E",X"E5",X"E6",X"07",X"21",X"88",X"34",
		X"CD",X"52",X"21",X"4E",X"E1",X"3A",X"51",X"4C",X"47",X"AF",X"81",X"10",X"FD",X"32",X"59",X"4C",
		X"C9",X"E5",X"F5",X"CD",X"3D",X"33",X"F1",X"4F",X"CD",X"4D",X"33",X"E1",X"C9",X"7E",X"0F",X"0F",
		X"E6",X"3E",X"21",X"90",X"34",X"CD",X"52",X"21",X"5E",X"23",X"56",X"EB",X"C9",X"11",X"4B",X"4C",
		X"E6",X"03",X"C4",X"6A",X"33",X"11",X"46",X"4C",X"79",X"0F",X"0F",X"4F",X"E6",X"03",X"C4",X"6A",
		X"33",X"11",X"41",X"4C",X"79",X"0F",X"0F",X"E6",X"03",X"C8",X"E5",X"3D",X"28",X"09",X"C5",X"44",
		X"4D",X"09",X"3D",X"28",X"01",X"09",X"C1",X"EB",X"7B",X"D7",X"77",X"23",X"7A",X"77",X"23",X"7A",
		X"D7",X"77",X"23",X"36",X"00",X"E1",X"C9",X"21",X"59",X"4C",X"7E",X"35",X"B7",X"E5",X"CC",X"D4",
		X"32",X"E1",X"2B",X"7E",X"34",X"2B",X"B7",X"20",X"0A",X"E5",X"CB",X"BE",X"2B",X"CB",X"BE",X"2B",
		X"CB",X"BE",X"E1",X"4F",X"7E",X"11",X"4F",X"4C",X"CD",X"BB",X"33",X"2B",X"7E",X"11",X"4A",X"4C",
		X"CD",X"BB",X"33",X"2B",X"7E",X"11",X"45",X"4C",X"C3",X"BB",X"33",X"87",X"C8",X"D8",X"E5",X"21",
		X"47",X"34",X"E6",X"1E",X"CD",X"52",X"21",X"7E",X"23",X"66",X"6F",X"79",X"0F",X"E6",X"7F",X"CD",
		X"52",X"21",X"7E",X"B7",X"E1",X"28",X"07",X"CB",X"41",X"20",X"01",X"D7",X"12",X"C9",X"CB",X"FE",
		X"C9",X"CB",X"BE",X"21",X"D0",X"34",X"11",X"6C",X"4C",X"C3",X"1F",X"34",X"CB",X"BE",X"11",X"60",
		X"4C",X"21",X"DC",X"34",X"C3",X"1F",X"34",X"CB",X"BE",X"11",X"6C",X"4C",X"21",X"E8",X"34",X"C3",
		X"1F",X"34",X"CB",X"BE",X"21",X"F4",X"34",X"CB",X"57",X"28",X"03",X"21",X"0C",X"35",X"11",X"60",
		X"4C",X"C3",X"1F",X"34",X"CB",X"BE",X"21",X"00",X"35",X"11",X"F0",X"4C",X"C3",X"1F",X"34",X"CB",
		X"7F",X"28",X"07",X"D5",X"01",X"0C",X"00",X"ED",X"B0",X"D1",X"D5",X"CD",X"38",X"34",X"CD",X"87",
		X"33",X"D1",X"CD",X"38",X"34",X"C3",X"E3",X"2D",X"21",X"50",X"4C",X"06",X"0C",X"1A",X"4E",X"77",
		X"79",X"12",X"23",X"13",X"10",X"F7",X"C9",X"00",X"00",X"59",X"34",X"62",X"34",X"6A",X"34",X"72",
		X"34",X"7C",X"34",X"7E",X"34",X"80",X"34",X"84",X"34",X"36",X"9C",X"EF",X"EB",X"98",X"76",X"66",
		X"55",X"00",X"13",X"57",X"99",X"75",X"54",X"33",X"22",X"00",X"7C",X"FF",X"EB",X"A8",X"77",X"65",
		X"54",X"00",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"00",X"55",X"00",X"FF",X"00",
		X"5C",X"5C",X"5C",X"00",X"12",X"23",X"34",X"00",X"01",X"02",X"04",X"06",X"08",X"0C",X"10",X"20",
		X"00",X"00",X"DC",X"09",X"89",X"0A",X"2B",X"0B",X"F3",X"0B",X"88",X"0C",X"46",X"0D",X"0C",X"0E",
		X"E6",X"0E",X"C9",X"0F",X"BA",X"10",X"B8",X"11",X"C6",X"12",X"E4",X"13",X"12",X"15",X"56",X"16",
		X"E7",X"17",X"10",X"19",X"8C",X"1A",X"21",X"1C",X"CC",X"1D",X"93",X"1F",X"74",X"21",X"70",X"23",
		X"8C",X"25",X"C7",X"27",X"25",X"2A",X"AC",X"2C",X"CF",X"2F",X"20",X"32",X"18",X"35",X"00",X"00",
		X"01",X"01",X"00",X"04",X"02",X"00",X"02",X"05",X"00",X"00",X"18",X"36",X"00",X"01",X"00",X"00",
		X"1C",X"04",X"04",X"00",X"00",X"00",X"40",X"36",X"01",X"01",X"00",X"0C",X"02",X"00",X"05",X"06",
		X"00",X"00",X"6B",X"36",X"01",X"01",X"00",X"0C",X"20",X"06",X"05",X"00",X"00",X"00",X"94",X"36",
		X"00",X"01",X"00",X"00",X"10",X"08",X"00",X"00",X"00",X"00",X"D4",X"36",X"01",X"01",X"00",X"08",
		X"20",X"06",X"06",X"00",X"00",X"00",X"1C",X"37",X"00",X"3E",X"00",X"32",X"4F",X"50",X"3E",X"01",
		X"32",X"4A",X"50",X"3E",X"02",X"32",X"45",X"50",X"F7",X"92",X"92",X"72",X"72",X"4C",X"4C",X"6C",
		X"AC",X"74",X"B4",X"92",X"92",X"72",X"72",X"4C",X"4C",X"6C",X"AC",X"74",X"B4",X"92",X"92",X"72",
		X"72",X"4C",X"4C",X"6A",X"AA",X"72",X"B2",X"34",X"34",X"72",X"B2",X"72",X"B2",X"24",X"24",X"74",
		X"A4",X"74",X"A4",X"92",X"92",X"72",X"72",X"24",X"24",X"74",X"A4",X"74",X"A4",X"92",X"92",X"72",
		X"72",X"24",X"24",X"74",X"A4",X"74",X"A4",X"92",X"92",X"72",X"72",X"24",X"24",X"72",X"A2",X"72",
		X"A2",X"34",X"34",X"72",X"A2",X"72",X"A2",X"4C",X"4C",X"6C",X"AC",X"74",X"B4",X"F9",X"F9",X"00",
		X"AF",X"21",X"5C",X"4C",X"77",X"23",X"77",X"23",X"77",X"23",X"36",X"81",X"CD",X"E0",X"2D",X"00",
		X"00",X"00",X"00",X"F7",X"F9",X"F9",X"00",X"3E",X"04",X"32",X"4F",X"50",X"3E",X"06",X"32",X"4A",
		X"50",X"F7",X"59",X"81",X"89",X"A9",X"59",X"81",X"89",X"A9",X"51",X"79",X"81",X"A1",X"51",X"79",
		X"81",X"A1",X"59",X"81",X"89",X"A9",X"59",X"81",X"89",X"A9",X"61",X"81",X"91",X"B1",X"61",X"81",
		X"91",X"B1",X"00",X"21",X"96",X"35",X"E5",X"C3",X"30",X"00",X"00",X"3E",X"06",X"32",X"45",X"50",
		X"3E",X"00",X"32",X"4A",X"50",X"F7",X"B3",X"A9",X"B3",X"C1",X"B4",X"FC",X"53",X"49",X"53",X"61",
		X"54",X"FC",X"B3",X"B1",X"FB",X"B1",X"C4",X"D4",X"DC",X"00",X"3E",X"01",X"32",X"51",X"4C",X"F7",
		X"18",X"20",X"28",X"30",X"38",X"40",X"48",X"50",X"58",X"60",X"68",X"70",X"78",X"80",X"88",X"90",
		X"98",X"A0",X"A8",X"B0",X"B8",X"C0",X"C8",X"D0",X"D8",X"E0",X"E8",X"F0",X"F8",X"00",X"3E",X"81",
		X"32",X"5C",X"4C",X"CD",X"E0",X"2D",X"F7",X"F9",X"00",X"3E",X"01",X"32",X"4A",X"50",X"3E",X"02",
		X"32",X"4F",X"50",X"F7",X"40",X"B8",X"58",X"B0",X"70",X"A8",X"58",X"A0",X"40",X"98",X"50",X"90",
		X"68",X"88",X"80",X"80",X"68",X"78",X"50",X"70",X"00",X"21",X"5E",X"4C",X"36",X"00",X"F7",X"F9",
		X"00",X"3E",X"04",X"32",X"45",X"50",X"3E",X"07",X"32",X"4A",X"50",X"F7",X"80",X"90",X"A0",X"B0",
		X"C0",X"D0",X"E0",X"F0",X"E0",X"D0",X"C0",X"B0",X"A0",X"90",X"80",X"90",X"80",X"90",X"A0",X"B0",
		X"C0",X"D0",X"E0",X"00",X"21",X"40",X"36",X"E5",X"C3",X"30",X"00",X"00",X"3E",X"01",X"32",X"4A",
		X"50",X"3E",X"03",X"32",X"4F",X"50",X"F7",X"08",X"A8",X"18",X"98",X"28",X"88",X"38",X"78",X"48",
		X"68",X"58",X"58",X"68",X"48",X"78",X"38",X"88",X"28",X"98",X"18",X"A8",X"08",X"00",X"21",X"6B",
		X"36",X"E5",X"F7",X"F9",X"00",X"3E",X"01",X"32",X"45",X"50",X"3E",X"03",X"32",X"4A",X"50",X"F7",
		X"40",X"B8",X"58",X"B0",X"78",X"A8",X"D8",X"A0",X"40",X"98",X"00",X"3E",X"07",X"32",X"45",X"50",
		X"3E",X"04",X"32",X"4A",X"50",X"F7",X"50",X"90",X"68",X"88",X"80",X"80",X"68",X"78",X"50",X"70",
		X"68",X"68",X"80",X"60",X"98",X"58",X"A8",X"50",X"98",X"48",X"80",X"40",X"00",X"21",X"5D",X"4C",
		X"36",X"00",X"F7",X"F9",X"00",X"3E",X"07",X"32",X"45",X"50",X"F7",X"62",X"39",X"39",X"62",X"39",
		X"39",X"99",X"99",X"89",X"89",X"7C",X"62",X"39",X"39",X"61",X"39",X"39",X"99",X"99",X"89",X"89",
		X"7C",X"00",X"3E",X"07",X"32",X"45",X"50",X"F7",X"61",X"61",X"71",X"71",X"79",X"79",X"89",X"89",
		X"79",X"79",X"71",X"71",X"61",X"61",X"72",X"61",X"61",X"71",X"71",X"79",X"79",X"89",X"89",X"79",
		X"79",X"71",X"71",X"64",X"00",X"21",X"D4",X"36",X"E5",X"C3",X"30",X"00",X"00",X"3E",X"01",X"32",
		X"45",X"50",X"3E",X"01",X"32",X"4A",X"50",X"F7",X"81",X"79",X"91",X"69",X"A1",X"59",X"B1",X"49",
		X"C1",X"39",X"B1",X"49",X"A1",X"59",X"91",X"69",X"81",X"79",X"00",X"21",X"78",X"4C",X"34",X"7E",
		X"FE",X"0A",X"28",X"07",X"21",X"1C",X"37",X"E5",X"C3",X"30",X"00",X"36",X"00",X"21",X"5D",X"4C",
		X"36",X"00",X"F7",X"09",X"97",X"F9",X"B4",X"35",X"11",X"00",X"C6",X"12",X"F9",X"E0",X"00",X"00",
		X"11",X"00",X"CD",X"12",X"B0",X"CB",X"96",X"00",X"52",X"37",X"11",X"00",X"DE",X"12",X"B0",X"CB",
		X"96",X"50",X"64",X"37",X"11",X"00",X"DF",X"12",X"F9",X"DE",X"00",X"00",X"11",X"00",X"E9",X"12",
		X"F9",X"DC",X"06",X"40",X"11",X"00",X"F2",X"12",X"F9",X"DC",X"0C",X"80",X"11",X"00",X"FF",X"12",
		X"F9",X"E1",X"00",X"00",X"11",X"00",X"05",X"13",X"F9",X"DD",X"00",X"00",X"11",X"00",X"07",X"13",
		X"F9",X"DA",X"00",X"00",X"11",X"00",X"0A",X"13",X"F9",X"DB",X"00",X"00",X"11",X"00",X"12",X"13",
		X"B0",X"CB",X"98",X"21",X"6E",X"37",X"11",X"00",X"1F",X"13",X"BF",X"58",X"8D",X"35",X"CB",X"32",
		X"11",X"00",X"27",X"13",X"F9",X"DB",X"00",X"00",X"11",X"00",X"2A",X"13",X"F9",X"DA",X"00",X"00",
		X"11",X"00",X"44",X"13",X"BF",X"56",X"A4",X"9A",X"9C",X"34",X"11",X"00",X"49",X"13",X"F9",X"DC",
		X"00",X"00",X"11",X"00",X"4E",X"13",X"F9",X"DA",X"00",X"00",X"11",X"00",X"5A",X"13",X"F9",X"DB",
		X"00",X"00",X"11",X"00",X"5B",X"13",X"BF",X"56",X"59",X"56",X"D4",X"37",X"11",X"00",X"5F",X"0D",
		X"C9",X"36",X"81",X"C3",X"E9",X"3E",X"C3",X"A8",X"2B",X"CD",X"3B",X"39",X"3A",X"C1",X"4F",X"B7",
		X"CA",X"0A",X"39",X"CB",X"67",X"21",X"E4",X"4F",X"20",X"1B",X"CB",X"77",X"7E",X"20",X"10",X"FE",
		X"50",X"28",X"2E",X"FE",X"18",X"CA",X"B2",X"38",X"FE",X"C0",X"28",X"45",X"C3",X"E8",X"38",X"B7",
		X"28",X"4B",X"C3",X"E8",X"38",X"CB",X"6F",X"7E",X"20",X"0C",X"FE",X"C0",X"28",X"47",X"FE",X"58",
		X"CA",X"DC",X"38",X"C3",X"E8",X"38",X"FE",X"02",X"30",X"F9",X"3E",X"0F",X"32",X"C0",X"4F",X"18",
		X"F2",X"2E",X"D8",X"36",X"22",X"23",X"23",X"36",X"22",X"2E",X"E8",X"36",X"10",X"23",X"36",X"60",
		X"23",X"36",X"01",X"23",X"36",X"60",X"3E",X"80",X"32",X"92",X"4C",X"32",X"94",X"4C",X"C3",X"E8",
		X"38",X"2E",X"D4",X"36",X"44",X"21",X"C1",X"4F",X"CB",X"F6",X"C3",X"E8",X"38",X"21",X"C1",X"4F",
		X"CB",X"E6",X"C3",X"E8",X"38",X"2E",X"D8",X"36",X"44",X"23",X"23",X"36",X"44",X"2E",X"C8",X"36",
		X"E0",X"23",X"36",X"07",X"23",X"36",X"E0",X"23",X"36",X"05",X"3E",X"40",X"32",X"32",X"42",X"32",
		X"52",X"42",X"E5",X"21",X"F7",X"41",X"06",X"07",X"11",X"20",X"00",X"77",X"19",X"10",X"FC",X"E1",
		X"18",X"A7",X"21",X"CC",X"4F",X"36",X"C0",X"23",X"36",X"07",X"2E",X"EC",X"36",X"00",X"23",X"36",
		X"60",X"2E",X"DC",X"36",X"44",X"3E",X"0D",X"32",X"96",X"4C",X"21",X"06",X"4E",X"36",X"00",X"23",
		X"36",X"01",X"23",X"3E",X"FF",X"77",X"32",X"10",X"4E",X"C3",X"E8",X"38",X"2E",X"D4",X"36",X"22",
		X"21",X"C1",X"4F",X"CB",X"EE",X"CD",X"94",X"3A",X"CD",X"55",X"2D",X"CD",X"C6",X"15",X"CD",X"40",
		X"26",X"CD",X"1D",X"0A",X"CD",X"81",X"09",X"CD",X"6A",X"11",X"CD",X"0A",X"20",X"CD",X"27",X"13",
		X"CD",X"E4",X"2A",X"CD",X"97",X"2C",X"CD",X"ED",X"2C",X"C9",X"21",X"E4",X"4F",X"36",X"10",X"23",
		X"36",X"60",X"21",X"33",X"39",X"11",X"C4",X"4F",X"01",X"08",X"00",X"ED",X"B0",X"21",X"D4",X"4F",
		X"36",X"22",X"3E",X"01",X"32",X"C1",X"4F",X"3E",X"0F",X"32",X"CE",X"4F",X"21",X"05",X"00",X"22",
		X"0E",X"4E",X"C9",X"F8",X"01",X"00",X"00",X"E0",X"07",X"E0",X"05",X"3A",X"C8",X"4F",X"CB",X"5F",
		X"28",X"04",X"AF",X"32",X"92",X"4C",X"3A",X"CA",X"4F",X"CB",X"5F",X"C8",X"AF",X"32",X"94",X"4C",
		X"C9",X"21",X"C1",X"4F",X"7E",X"34",X"FE",X"80",X"D8",X"21",X"C0",X"4F",X"36",X"1F",X"C9",X"7E",
		X"FE",X"04",X"D0",X"3A",X"5C",X"4C",X"FE",X"03",X"C0",X"36",X"05",X"C9",X"3E",X"19",X"21",X"2A",
		X"46",X"11",X"1D",X"00",X"0E",X"04",X"C3",X"A7",X"28",X"3E",X"19",X"21",X"6A",X"45",X"11",X"1D",
		X"00",X"0E",X"04",X"C3",X"A7",X"28",X"11",X"C8",X"4F",X"21",X"EE",X"4F",X"7E",X"B7",X"28",X"0E",
		X"35",X"20",X"07",X"06",X"A0",X"CD",X"AE",X"39",X"18",X"04",X"AF",X"32",X"92",X"4C",X"23",X"13",
		X"13",X"7E",X"B7",X"C8",X"35",X"06",X"70",X"28",X"05",X"AF",X"32",X"94",X"4C",X"C9",X"D5",X"E5",
		X"23",X"23",X"36",X"00",X"E1",X"EB",X"36",X"48",X"23",X"36",X"09",X"7D",X"C6",X"1F",X"6F",X"70",
		X"23",X"36",X"B0",X"7D",X"D6",X"31",X"6F",X"36",X"00",X"C6",X"20",X"6F",X"36",X"10",X"EB",X"E5",
		X"CD",X"29",X"10",X"E1",X"D1",X"3A",X"48",X"50",X"07",X"C9",X"3A",X"8D",X"50",X"E6",X"C0",X"C8",
		X"87",X"87",X"D8",X"00",X"00",X"21",X"12",X"4E",X"34",X"C9",X"3A",X"20",X"4C",X"E6",X"03",X"C8",
		X"3A",X"06",X"4E",X"32",X"9F",X"4C",X"C9",X"16",X"01",X"7D",X"1E",X"10",X"FE",X"05",X"C8",X"1E",
		X"14",X"FE",X"10",X"C8",X"1E",X"18",X"FE",X"20",X"20",X"06",X"7C",X"B7",X"C8",X"1E",X"38",X"C9",
		X"1E",X"1C",X"FE",X"40",X"20",X"06",X"7C",X"B7",X"C8",X"1E",X"3C",X"C9",X"1E",X"30",X"FE",X"80",
		X"C8",X"1E",X"34",X"FE",X"60",X"C8",X"1E",X"50",X"C9",X"1A",X"85",X"27",X"12",X"1B",X"1A",X"8C",
		X"27",X"12",X"1B",X"1A",X"CE",X"00",X"27",X"12",X"C9",X"7D",X"32",X"0C",X"4E",X"85",X"27",X"6F",
		X"7C",X"32",X"0B",X"4E",X"8C",X"27",X"67",X"3E",X"FF",X"32",X"0D",X"4E",X"D0",X"21",X"99",X"99",
		X"C9",X"7D",X"D6",X"30",X"6F",X"7B",X"D6",X"30",X"5F",X"1A",X"AE",X"E6",X"80",X"C8",X"C3",X"7E",
		X"3A",X"E5",X"D5",X"CD",X"76",X"3A",X"D1",X"E1",X"3E",X"7F",X"20",X"07",X"CD",X"9A",X"2B",X"4F",
		X"C3",X"9A",X"2B",X"23",X"23",X"C9",X"7D",X"D6",X"10",X"6F",X"7B",X"D6",X"10",X"5F",X"1A",X"B6",
		X"E6",X"0F",X"FE",X"09",X"C8",X"FE",X"06",X"C8",X"FE",X"01",X"C8",X"FE",X"02",X"C8",X"FE",X"04",
		X"C8",X"FE",X"08",X"C9",X"3A",X"81",X"4C",X"FE",X"20",X"D8",X"E5",X"21",X"BC",X"42",X"11",X"20",
		X"00",X"06",X"05",X"AF",X"86",X"19",X"10",X"FC",X"FE",X"65",X"E1",X"C8",X"3E",X"01",X"32",X"01",
		X"4C",X"32",X"20",X"4C",X"C9",X"3E",X"01",X"32",X"04",X"50",X"21",X"D0",X"4C",X"34",X"7E",X"FE",
		X"3C",X"D8",X"36",X"00",X"23",X"34",X"7E",X"FE",X"1E",X"D8",X"AF",X"77",X"32",X"04",X"50",X"C9",
		X"3A",X"D1",X"4C",X"FE",X"07",X"C8",X"FE",X"0B",X"C8",X"87",X"E6",X"7E",X"21",X"BD",X"0E",X"CD",
		X"52",X"21",X"3A",X"C0",X"50",X"E6",X"00",X"00",X"C9",X"23",X"3A",X"80",X"50",X"86",X"C0",X"B0",
		X"C9",X"21",X"9D",X"4C",X"7E",X"B7",X"C8",X"35",X"C0",X"23",X"36",X"00",X"C9",X"E5",X"D5",X"7D",
		X"C6",X"10",X"6F",X"7E",X"FE",X"88",X"28",X"06",X"56",X"21",X"32",X"3B",X"18",X"06",X"23",X"56",
		X"2B",X"21",X"3E",X"3B",X"CD",X"1D",X"3B",X"D1",X"E1",X"D4",X"C5",X"1A",X"C9",X"3A",X"9E",X"4C",
		X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"E6",X"0E",X"CD",X"52",X"21",X"7A",X"BE",X"D8",X"23",X"BE",
		X"3F",X"C9",X"18",X"FF",X"20",X"F8",X"28",X"F0",X"30",X"E8",X"40",X"D8",X"50",X"C8",X"20",X"FF",
		X"30",X"FF",X"40",X"FF",X"50",X"F8",X"60",X"F0",X"6C",X"E8",X"3A",X"83",X"4C",X"E6",X"7F",X"FE",
		X"75",X"C0",X"ED",X"5F",X"85",X"83",X"E6",X"03",X"CD",X"8F",X"3B",X"1A",X"CB",X"7F",X"C0",X"E6",
		X"7F",X"FE",X"10",X"D0",X"E5",X"CD",X"A7",X"3B",X"E1",X"C0",X"E5",X"7C",X"C6",X"04",X"67",X"CD",
		X"B4",X"3B",X"E1",X"C0",X"D5",X"E5",X"CD",X"D7",X"3B",X"D1",X"E1",X"34",X"CB",X"FE",X"EB",X"06",
		X"BE",X"70",X"23",X"04",X"70",X"04",X"CD",X"50",X"21",X"2B",X"70",X"04",X"23",X"70",X"C9",X"11",
		X"1E",X"4E",X"21",X"A8",X"42",X"C8",X"13",X"21",X"28",X"41",X"3D",X"C8",X"13",X"21",X"B1",X"42",
		X"3D",X"C8",X"13",X"21",X"31",X"41",X"C9",X"7E",X"23",X"A6",X"F5",X"CD",X"50",X"21",X"F1",X"A6",
		X"2B",X"A6",X"3C",X"C9",X"7E",X"E6",X"1F",X"FE",X"02",X"28",X"07",X"FE",X"04",X"28",X"03",X"FE",
		X"06",X"C0",X"47",X"23",X"7E",X"E6",X"1F",X"B8",X"C0",X"CD",X"50",X"21",X"7E",X"E6",X"1F",X"B8",
		X"C0",X"2B",X"7E",X"E6",X"1F",X"B8",X"C9",X"CD",X"E5",X"3B",X"21",X"1E",X"4E",X"06",X"04",X"CB",
		X"BE",X"23",X"10",X"FB",X"C9",X"11",X"1E",X"4E",X"21",X"A8",X"42",X"CD",X"FD",X"3B",X"21",X"28",
		X"41",X"CD",X"FD",X"3B",X"21",X"B1",X"42",X"CD",X"FD",X"3B",X"21",X"31",X"41",X"1A",X"13",X"87",
		X"D0",X"06",X"FF",X"70",X"23",X"70",X"CD",X"50",X"21",X"70",X"2B",X"70",X"C9",X"7A",X"D6",X"BE",
		X"C8",X"3D",X"C8",X"3D",X"C8",X"3D",X"C9",X"2A",X"E4",X"4F",X"7D",X"FE",X"B8",X"28",X"1B",X"FE",
		X"58",X"C0",X"7C",X"FE",X"C0",X"28",X"0B",X"FE",X"78",X"C0",X"21",X"31",X"41",X"11",X"21",X"4E",
		X"18",X"1E",X"21",X"28",X"41",X"11",X"1F",X"4E",X"18",X"16",X"7C",X"FE",X"C0",X"28",X"0B",X"FE",
		X"78",X"C0",X"21",X"B1",X"42",X"11",X"20",X"4E",X"18",X"06",X"21",X"A8",X"42",X"11",X"1E",X"4E",
		X"1A",X"07",X"D0",X"EB",X"CB",X"BE",X"EB",X"CD",X"01",X"3C",X"21",X"88",X"18",X"22",X"E4",X"4F",
		X"C9",X"11",X"1E",X"4E",X"21",X"A8",X"42",X"CD",X"79",X"3C",X"21",X"28",X"41",X"CD",X"79",X"3C",
		X"21",X"B1",X"42",X"CD",X"79",X"3C",X"21",X"31",X"41",X"1A",X"13",X"87",X"D0",X"C3",X"7F",X"3B",
		X"3A",X"AE",X"4C",X"B7",X"28",X"06",X"CD",X"C4",X"1D",X"C3",X"86",X"03",X"3A",X"AC",X"4C",X"07",
		X"38",X"0D",X"21",X"AF",X"4C",X"35",X"20",X"04",X"AF",X"32",X"AC",X"4C",X"C3",X"86",X"03",X"3E",
		X"01",X"32",X"AC",X"4C",X"3E",X"FF",X"32",X"AF",X"4C",X"21",X"E0",X"4F",X"06",X"20",X"36",X"00",
		X"23",X"10",X"FB",X"3E",X"03",X"CD",X"5B",X"2E",X"CD",X"50",X"0D",X"CD",X"38",X"22",X"CD",X"DD",
		X"3C",X"CD",X"C7",X"3C",X"C3",X"86",X"03",X"3E",X"01",X"01",X"E0",X"FF",X"11",X"40",X"4E",X"21",
		X"CB",X"42",X"F5",X"CD",X"0F",X"3D",X"F1",X"3C",X"FE",X"06",X"20",X"F6",X"C9",X"CD",X"DF",X"0C",
		X"CD",X"02",X"0D",X"CD",X"80",X"28",X"0F",X"08",X"41",X"53",X"52",X"45",X"59",X"41",X"4C",X"50",
		X"40",X"54",X"55",X"4F",X"40",X"52",X"41",X"46",X"21",X"08",X"45",X"06",X"0F",X"36",X"01",X"CD",
		X"50",X"21",X"10",X"F9",X"21",X"CB",X"46",X"06",X"0C",X"36",X"05",X"23",X"10",X"FB",X"C9",X"E5",
		X"77",X"09",X"09",X"3E",X"03",X"08",X"1A",X"77",X"13",X"09",X"08",X"3D",X"20",X"F7",X"09",X"CD",
		X"26",X"3D",X"E1",X"23",X"23",X"C9",X"3E",X"03",X"08",X"1A",X"D7",X"E6",X"0F",X"20",X"15",X"09",
		X"1A",X"E6",X"0F",X"20",X"14",X"09",X"13",X"08",X"3D",X"20",X"ED",X"08",X"36",X"00",X"C9",X"08",
		X"1A",X"D7",X"E6",X"0F",X"77",X"09",X"1A",X"E6",X"0F",X"77",X"09",X"13",X"08",X"3D",X"20",X"EF",
		X"18",X"E9",X"78",X"32",X"68",X"4E",X"B7",X"20",X"05",X"7E",X"E6",X"7D",X"77",X"C9",X"CB",X"7E",
		X"20",X"2D",X"CD",X"F9",X"0E",X"3A",X"AF",X"4C",X"B7",X"C0",X"21",X"AE",X"4C",X"18",X"EA",X"79",
		X"32",X"68",X"4E",X"B7",X"20",X"08",X"7E",X"E6",X"86",X"77",X"CD",X"D7",X"2D",X"C9",X"CB",X"76",
		X"20",X"2D",X"CD",X"F9",X"0E",X"3A",X"AF",X"4C",X"B7",X"C0",X"21",X"AE",X"4C",X"18",X"E7",X"CB",
		X"BE",X"F5",X"CD",X"D7",X"2D",X"F1",X"CD",X"D8",X"3D",X"CD",X"6B",X"0F",X"36",X"41",X"AF",X"12",
		X"CD",X"80",X"28",X"07",X"84",X"41",X"01",X"52",X"45",X"59",X"41",X"4C",X"50",X"18",X"23",X"CB",
		X"B6",X"F5",X"3A",X"00",X"50",X"CB",X"67",X"C4",X"DA",X"2D",X"F1",X"CD",X"D8",X"3D",X"CD",X"6B",
		X"0F",X"36",X"41",X"AF",X"12",X"CD",X"80",X"28",X"07",X"84",X"41",X"02",X"52",X"45",X"59",X"41",
		X"4C",X"50",X"3E",X"40",X"32",X"AF",X"4C",X"C9",X"F5",X"3E",X"03",X"CD",X"5B",X"2E",X"CD",X"50",
		X"0D",X"CD",X"38",X"22",X"CD",X"E3",X"3C",X"CD",X"C7",X"3C",X"CD",X"F1",X"3D",X"F1",X"C3",X"9B",
		X"3E",X"CD",X"80",X"28",X"15",X"C6",X"40",X"53",X"4C",X"41",X"49",X"54",X"49",X"4E",X"49",X"40",
		X"52",X"55",X"4F",X"59",X"40",X"4E",X"47",X"49",X"53",X"40",X"4F",X"54",X"21",X"C6",X"44",X"06",
		X"15",X"36",X"05",X"CD",X"50",X"21",X"10",X"F9",X"CD",X"80",X"28",X"13",X"D5",X"40",X"48",X"54",
		X"49",X"57",X"40",X"4C",X"41",X"49",X"54",X"49",X"4E",X"49",X"40",X"54",X"43",X"45",X"4C",X"45",
		X"53",X"CD",X"80",X"28",X"10",X"16",X"41",X"54",X"46",X"45",X"4C",X"40",X"40",X"44",X"4E",X"41",
		X"40",X"40",X"54",X"48",X"47",X"49",X"52",X"CD",X"80",X"28",X"0D",X"78",X"41",X"4E",X"57",X"4F",
		X"44",X"40",X"48",X"54",X"49",X"57",X"40",X"42",X"55",X"52",X"CD",X"80",X"28",X"0D",X"79",X"41",
		X"50",X"55",X"40",X"48",X"54",X"49",X"57",X"40",X"45",X"54",X"49",X"52",X"57",X"21",X"D5",X"44",
		X"0E",X"05",X"E5",X"06",X"13",X"36",X"05",X"CD",X"50",X"21",X"10",X"F9",X"E1",X"23",X"0D",X"20",
		X"F1",X"CD",X"80",X"28",X"07",X"DB",X"41",X"00",X"04",X"40",X"45",X"4D",X"49",X"54",X"21",X"84",
		X"45",X"06",X"07",X"36",X"07",X"CD",X"50",X"21",X"10",X"F9",X"C9",X"21",X"0B",X"45",X"D6",X"05",
		X"ED",X"44",X"87",X"CD",X"52",X"21",X"06",X"0F",X"36",X"01",X"CD",X"50",X"21",X"10",X"F9",X"C9",
		X"3A",X"83",X"4C",X"E6",X"3F",X"FE",X"17",X"C0",X"21",X"AF",X"4C",X"7E",X"D6",X"01",X"27",X"77",
		X"D7",X"E6",X"0F",X"20",X"02",X"3E",X"40",X"32",X"FB",X"41",X"7E",X"E6",X"0F",X"32",X"DB",X"41",
		X"C9",X"00",X"19",X"19",X"B8",X"29",X"B3",X"B0",X"C2",X"3E",X"11",X"00",X"1C",X"19",X"B8",X"29",
		X"3A",X"80",X"50",X"CB",X"6F",X"C8",X"C3",X"A8",X"2B",X"3A",X"80",X"50",X"E6",X"3F",X"C0",X"3E",
		X"03",X"CD",X"5B",X"2E",X"3E",X"40",X"CD",X"65",X"2E",X"CD",X"80",X"28",X"06",X"89",X"40",X"57",
		X"53",X"40",X"50",X"49",X"44",X"0E",X"00",X"3A",X"80",X"50",X"E6",X"3F",X"47",X"3A",X"80",X"50",
		X"A8",X"E6",X"3F",X"B1",X"FE",X"3F",X"28",X"06",X"4F",X"32",X"C0",X"50",X"18",X"EF",X"3E",X"40",
		X"CD",X"65",X"2E",X"21",X"D0",X"4C",X"36",X"00",X"23",X"10",X"FB",X"CD",X"80",X"28",X"0A",X"83",
		X"40",X"4B",X"48",X"43",X"40",X"4D",X"55",X"54",X"53",X"55",X"43",X"3E",X"01",X"32",X"04",X"50",
		X"32",X"07",X"50",X"0E",X"04",X"32",X"C0",X"50",X"10",X"FB",X"0D",X"20",X"F8",X"AF",X"32",X"04",
		X"50",X"21",X"D0",X"4C",X"77",X"23",X"77",X"23",X"77",X"21",X"D0",X"4C",X"7E",X"2F",X"32",X"07",
		X"50",X"32",X"C0",X"50",X"2F",X"34",X"FE",X"78",X"20",X"08",X"36",X"00",X"23",X"34",X"7E",X"FE",
		X"1E",X"C8",X"06",X"00",X"10",X"FE",X"3A",X"D0",X"4C",X"FE",X"10",X"38",X"DC",X"FE",X"6E",X"30",
		X"D8",X"CD",X"D0",X"3A",X"28",X"D3",X"CD",X"80",X"28",X"05",X"85",X"40",X"52",X"52",X"4F",X"52",
		X"45",X"32",X"C0",X"50",X"18",X"FB",X"CD",X"80",X"28",X"05",X"85",X"40",X"4B",X"4F",X"40",X"40",
		X"40",X"18",X"EE",X"00",X"2B",X"C9",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"FE",X"0A",X"38",
		X"02",X"C6",X"37",X"77",X"79",X"2B",X"E6",X"0F",X"FE",X"0A",X"38",X"02",X"C6",X"37",X"77",X"2B",
		X"C9",X"3C",X"8A",X"20",X"B6",X"3F",X"11",X"00",X"CD",X"80",X"3F",X"F5",X"F3",X"3A",X"00",X"50",
		X"CB",X"67",X"32",X"C0",X"50",X"28",X"F6",X"3A",X"00",X"50",X"CB",X"67",X"32",X"C0",X"50",X"20",
		X"F6",X"E5",X"21",X"00",X"50",X"36",X"00",X"36",X"01",X"E1",X"F1",X"FB",X"C9",X"3F",X"11",X"00",
		X"D2",X"1A",X"F9",X"DA",X"00",X"00",X"11",X"00",X"DC",X"1A",X"B8",X"29",X"BF",X"03",X"DE",X"A4");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
